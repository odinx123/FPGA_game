// 四倍小
module menu_img_160(clk, rst, X, Y, mapR, mapG, mapB);

	parameter xbit = 10, ybit = 9;
	input clk, rst;
	input [xbit-1:0] X;
	input [ybit-1:0] Y;
	output [7:0] mapR, mapG, mapB;
	reg [7:0] mapR, mapG, mapB;

	always @(posedge clk, negedge rst) begin
		if(!rst) begin
			mapR <= 8'd255;
			mapG <= 8'd255;
			mapB <= 8'd255;
		end
		else begin
			case(Y)
				`ybit'd0: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd209, 8'd222, 8'd254};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd210, 8'd222, 8'd254};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd210, 8'd222, 8'd253};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd209, 8'd222, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd211, 8'd221, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd211, 8'd221, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd254};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd253};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd212, 8'd221, 8'd249};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd211, 8'd221, 8'd248};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd212, 8'd221, 8'd250};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd212, 8'd221, 8'd250};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd214, 8'd223, 8'd252};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd214, 8'd223, 8'd252};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd252};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd250};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd249};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd253};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd213, 8'd223, 8'd250};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd213, 8'd222, 8'd251};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd213, 8'd222, 8'd251};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd249};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd213, 8'd225, 8'd250};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd213, 8'd225, 8'd250};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd213, 8'd225, 8'd250};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd212, 8'd221, 8'd252};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd251};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd211, 8'd223, 8'd251};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd211, 8'd223, 8'd251};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd211, 8'd223, 8'd251};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd252};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd253};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd253};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd211, 8'd221, 8'd255};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd211, 8'd221, 8'd255};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd211, 8'd221, 8'd255};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd255};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd254};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd254};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
					endcase
				end
				`ybit'd1: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd208, 8'd222, 8'd254};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd210, 8'd222, 8'd254};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd209, 8'd221, 8'd253};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd208, 8'd221, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd254};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd254};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd250};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd209, 8'd217, 8'd252};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd249};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd249};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd213, 8'd222, 8'd250};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd213, 8'd222, 8'd251};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd252};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd251};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd249};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd253};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd252};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd252};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd252};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd206, 8'd220, 8'd251};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd253};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd253};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd253};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd253};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd250};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd248};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd249};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd251};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd212, 8'd222, 8'd252};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd251};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd222, 8'd254};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd253};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd253};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd254};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd254};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd253};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd252};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd252};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd252};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd252};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd253};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd255};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd254};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd254};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd255};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
					endcase
				end
				`ybit'd2: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd208, 8'd217, 8'd252};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd252};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd252};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd253};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd209, 8'd219, 8'd253};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd250};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd253};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd253};
					endcase
				end
				`ybit'd3: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd251};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd247};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd240};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd241};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd246};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd251};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd251};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd251};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd250};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd252};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd252};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd252};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd251};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd251};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd251};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd251};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd252};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd250};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd250};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd250};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd250};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd250};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd250};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd250};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd207, 8'd217, 8'd250};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd206, 8'd218, 8'd250};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd250};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd251};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd252};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd206, 8'd218, 8'd250};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd251};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd252};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd251};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd252};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd250};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd251};
					endcase
				end
				`ybit'd4: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd206, 8'd218, 8'd245};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd202, 8'd214, 8'd239};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd196, 8'd209, 8'd229};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd196, 8'd209, 8'd228};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd202, 8'd214, 8'd240};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd247};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd249};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd250};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd250};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd249};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd250};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd249};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd250};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd250};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd205, 8'd215, 8'd250};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd205, 8'd215, 8'd250};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd205, 8'd215, 8'd250};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd203, 8'd216, 8'd250};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd251};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd251};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd251};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd250};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd249};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd206, 8'd219, 8'd251};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd206, 8'd219, 8'd251};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd206, 8'd219, 8'd251};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd251};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd250};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
					endcase
				end
				`ybit'd5: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd245};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd244};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd243};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd241};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd242};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd243};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd243};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd249};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd249};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd249};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd251};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd210, 8'd221, 8'd249};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd249};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd244};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd200, 8'd212, 8'd237};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd228};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd213};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd211};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd226};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd250};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd249};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd249};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd249};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd249};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd249};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd204, 8'd216, 8'd249};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd207, 8'd219, 8'd249};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd249};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd249};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd249};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd249};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
					endcase
				end
				`ybit'd6: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd248};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd201, 8'd213, 8'd239};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd231};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd194, 8'd206, 8'd227};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd194, 8'd207, 8'd228};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd194, 8'd206, 8'd227};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd195, 8'd208, 8'd227};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd228};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd197, 8'd210, 8'd231};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd201, 8'd213, 8'd236};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd248};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd248};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd248};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd247};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd246};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd246};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd247};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd241};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd234};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd189, 8'd202, 8'd220};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd184, 8'd197, 8'd207};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd176, 8'd189, 8'd198};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd175, 8'd188, 8'd196};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd212};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd232};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd209, 8'd220, 8'd250};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd247};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd248};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd203, 8'd216, 8'd248};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd203, 8'd216, 8'd248};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd203, 8'd216, 8'd248};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd203, 8'd216, 8'd248};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd203, 8'd216, 8'd248};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd204, 8'd217, 8'd249};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd205, 8'd218, 8'd250};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd249};
					endcase
				end
				`ybit'd7: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd234};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd189, 8'd200, 8'd220};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd181, 8'd193, 8'd208};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd180, 8'd192, 8'd206};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd182, 8'd194, 8'd207};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd181, 8'd195, 8'd203};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd181, 8'd195, 8'd203};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd213};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd194, 8'd206, 8'd228};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd201, 8'd213, 8'd238};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd241};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd242};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd243};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd201, 8'd213, 8'd238};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd232};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd198, 8'd208, 8'd233};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd199, 8'd211, 8'd231};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd200, 8'd212, 8'd239};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd200, 8'd212, 8'd239};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd197, 8'd208, 8'd230};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd215};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd179, 8'd191, 8'd200};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd173, 8'd183, 8'd189};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd167, 8'd178, 8'd182};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd167, 8'd178, 8'd180};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd179, 8'd189, 8'd198};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd227};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd240};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd245};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd245};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd246};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd246};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd246};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd246};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd206, 8'd216, 8'd246};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd248};
					endcase
				end
				`ybit'd8: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd238};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd193, 8'd206, 8'd224};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd181, 8'd193, 8'd208};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd172, 8'd180, 8'd187};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd167, 8'd175, 8'd180};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd165, 8'd179, 8'd180};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd165, 8'd181, 8'd180};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd165, 8'd181, 8'd180};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd170, 8'd185, 8'd189};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd182, 8'd196, 8'd207};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd193, 8'd205, 8'd224};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd234};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd200, 8'd213, 8'd238};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd240};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd196, 8'd208, 8'd236};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd196, 8'd208, 8'd230};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd196, 8'd208, 8'd230};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd234};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd199, 8'd211, 8'd236};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd199, 8'd211, 8'd235};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd229};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd229};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd229};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd232};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd235};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd235};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd200, 8'd213, 8'd238};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd201, 8'd213, 8'd238};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd194, 8'd207, 8'd225};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd199, 8'd210};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd210};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd187, 8'd200, 8'd215};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd190, 8'd202, 8'd224};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd189, 8'd202, 8'd223};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd208};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd175, 8'd189, 8'd193};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd165, 8'd179, 8'd177};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd161, 8'd174, 8'd170};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd161, 8'd173, 8'd171};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd163, 8'd174, 8'd176};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd173, 8'd184, 8'd193};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd188, 8'd200, 8'd218};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd229};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd231};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd232};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd231};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd232};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd198, 8'd211, 8'd235};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd200, 8'd212, 8'd237};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd240};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd244};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd246};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd246};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd205, 8'd217, 8'd247};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd206, 8'd217, 8'd247};
					endcase
				end
				`ybit'd9: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd243};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd200, 8'd211, 8'd239};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd196, 8'd208, 8'd230};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd172, 8'd186, 8'd195};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd161, 8'd172, 8'd175};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd154, 8'd166, 8'd163};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd152, 8'd167, 8'd158};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd153, 8'd168, 8'd159};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd153, 8'd169, 8'd159};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd159, 8'd174, 8'd172};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd169, 8'd183, 8'd188};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd179, 8'd193, 8'd203};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd214};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd190, 8'd203, 8'd224};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd235};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd200, 8'd212, 8'd238};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd195, 8'd206, 8'd230};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd187, 8'd200, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd183, 8'd196, 8'd210};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd183, 8'd195, 8'd213};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd213};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd189, 8'd201, 8'd222};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd191, 8'd203, 8'd223};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd187, 8'd200, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd214};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd214};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd215};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd215};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd187, 8'd200, 8'd215};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd191, 8'd203, 8'd225};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd196, 8'd208, 8'd235};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd201, 8'd211, 8'd241};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd243};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd243};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd242};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd196, 8'd208, 8'd235};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd212};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd173, 8'd186, 8'd193};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd170, 8'd183, 8'd190};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd173, 8'd186, 8'd195};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd178, 8'd190, 8'd200};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd176, 8'd188, 8'd198};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd170, 8'd183, 8'd189};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd162, 8'd175, 8'd173};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd156, 8'd169, 8'd160};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd157, 8'd166, 8'd159};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd157, 8'd168, 8'd166};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd160, 8'd169, 8'd172};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd173, 8'd181, 8'd191};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd183, 8'd195, 8'd210};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd215};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd213};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd189, 8'd197, 8'd212};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd187, 8'd197, 8'd208};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd210};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd215};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd219};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd193, 8'd205, 8'd224};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd230};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd235};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd199, 8'd209, 8'd234};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd201, 8'd209, 8'd239};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd202, 8'd211, 8'd236};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd200, 8'd214, 8'd239};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd204, 8'd212, 8'd243};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd244};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd244};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd202, 8'd215, 8'd242};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd243};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd202, 8'd215, 8'd243};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd201, 8'd214, 8'd243};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd205, 8'd214, 8'd245};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd244};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd244};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd244};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd245};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd242};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd246};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd245};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd202, 8'd215, 8'd245};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd202, 8'd215, 8'd245};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd245};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd202, 8'd215, 8'd245};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd246};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd245};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd202, 8'd216, 8'd245};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd202, 8'd216, 8'd245};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd202, 8'd215, 8'd245};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd245};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd205, 8'd213, 8'd249};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd245};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd205, 8'd214, 8'd244};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd246};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd205, 8'd214, 8'd244};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd203, 8'd215, 8'd244};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd204, 8'd215, 8'd245};
					endcase
				end
				`ybit'd10: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd241};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd197, 8'd208, 8'd236};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd189, 8'd202, 8'd223};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd177, 8'd191, 8'd203};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd165, 8'd179, 8'd184};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd155, 8'd167, 8'd165};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd148, 8'd161, 8'd152};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd145, 8'd161, 8'd148};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd145, 8'd161, 8'd147};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd145, 8'd161, 8'd148};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd150, 8'd165, 8'd157};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd157, 8'd172, 8'd166};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd164, 8'd179, 8'd179};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd170, 8'd185, 8'd190};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd178, 8'd192, 8'd204};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd190, 8'd202, 8'd223};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd195, 8'd207, 8'd233};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd189, 8'd202, 8'd221};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd175, 8'd189, 8'd199};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd168, 8'd183, 8'd186};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd168, 8'd182, 8'd183};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd169, 8'd184, 8'd188};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd174, 8'd188, 8'd200};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd179, 8'd191, 8'd207};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd202};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd175, 8'd189, 8'd196};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd172, 8'd187, 8'd193};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd171, 8'd186, 8'd191};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd171, 8'd185, 8'd191};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd171, 8'd185, 8'd190};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd175, 8'd189, 8'd201};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd215};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd194, 8'd206, 8'd229};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd238};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd242};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd200, 8'd211, 8'd239};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd193, 8'd206, 8'd227};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd178, 8'd192, 8'd200};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd163, 8'd177, 8'd179};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd158, 8'd173, 8'd169};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd160, 8'd174, 8'd175};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd163, 8'd177, 8'd178};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd161, 8'd176, 8'd172};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd155, 8'd170, 8'd165};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd151, 8'd164, 8'd156};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd149, 8'd162, 8'd149};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd151, 8'd161, 8'd151};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd61};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd146, 8'd139, 8'd135};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd144, 8'd136, 8'd136};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd100};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd177, 8'd186, 8'd192};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd173, 8'd184, 8'd185};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd100, 8'd102, 8'd104};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd141, 8'd136, 8'd135};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd146, 8'd137, 8'd136};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd80, 8'd77, 8'd77};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd81, 8'd78, 8'd78};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd145, 8'd139, 8'd135};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd137};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd121, 8'd122, 8'd126};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd150, 8'd140, 8'd139};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd145, 8'd137, 8'd134};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd155, 8'd145, 8'd143};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd223};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd99, 8'd101, 8'd107};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd145, 8'd136, 8'd134};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd145, 8'd135, 8'd134};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd100, 8'd101, 8'd108};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd139, 8'd130, 8'd130};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd145, 8'd135, 8'd136};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd145, 8'd136, 8'd136};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd148, 8'd137, 8'd136};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd147, 8'd136, 8'd135};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd143, 8'd137, 8'd132};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd152, 8'd147, 8'd141};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd63, 8'd60, 8'd58};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd133};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd133};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd143, 8'd137, 8'd134};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd143, 8'd136, 8'd133};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd146, 8'd139, 8'd136};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd148, 8'd137, 8'd135};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd128, 8'd128, 8'd128};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd145, 8'd137, 8'd134};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd129, 8'd123, 8'd119};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd144, 8'd137, 8'd134};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd135};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd133};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd143, 8'd137, 8'd133};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd99, 8'd102, 8'd107};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd150, 8'd143, 8'd147};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd146, 8'd137, 8'd133};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd147, 8'd138, 8'd135};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd145, 8'd136, 8'd134};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd146, 8'd135, 8'd133};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd145, 8'd136, 8'd134};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd151, 8'd143, 8'd142};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd14, 8'd16, 8'd20};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd144, 8'd135, 8'd133};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd146, 8'd137, 8'd134};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd145, 8'd137, 8'd134};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd128, 8'd119, 8'd117};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd147, 8'd137, 8'd135};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd148, 8'd140, 8'd131};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd124, 8'd124, 8'd131};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd149, 8'd138, 8'd134};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd148, 8'd137, 8'd136};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd146, 8'd135, 8'd133};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd131, 8'd121, 8'd119};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd144, 8'd135, 8'd132};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd73};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd204, 8'd212, 8'd243};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd244};
					endcase
				end
				`ybit'd11: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd199, 8'd213, 8'd240};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd195, 8'd208, 8'd235};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd185, 8'd200, 8'd219};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd174, 8'd188, 8'd197};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd160, 8'd175, 8'd175};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd150, 8'd165, 8'd161};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd145, 8'd161, 8'd150};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd142, 8'd158, 8'd148};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd140, 8'd156, 8'd145};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd141, 8'd157, 8'd147};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd143, 8'd160, 8'd150};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd150, 8'd162, 8'd155};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd152, 8'd167, 8'd161};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd158, 8'd172, 8'd172};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd169, 8'd183, 8'd188};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd182, 8'd195, 8'd211};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd191, 8'd203, 8'd224};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd184, 8'd197, 8'd212};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd168, 8'd183, 8'd185};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd155, 8'd172, 8'd165};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd154, 8'd169, 8'd161};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd153, 8'd168, 8'd163};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd160, 8'd174, 8'd176};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd166, 8'd180, 8'd185};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd169, 8'd183, 8'd187};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd166, 8'd180, 8'd182};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd161, 8'd175, 8'd178};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd159, 8'd173, 8'd170};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd155, 8'd169, 8'd166};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd156, 8'd171, 8'd166};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd161, 8'd175, 8'd177};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd172, 8'd184, 8'd193};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd184, 8'd195, 8'd213};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd193, 8'd205, 8'd226};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd197, 8'd209, 8'd236};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd199, 8'd211, 8'd238};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd236};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd190, 8'd203, 8'd222};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd173, 8'd188, 8'd194};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd160, 8'd173, 8'd173};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd156, 8'd167, 8'd166};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd155, 8'd167, 8'd163};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd156, 8'd168, 8'd164};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd153, 8'd166, 8'd155};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd149, 8'd162, 8'd149};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd146, 8'd160, 8'd147};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd144, 8'd158, 8'd145};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd150, 8'd156, 8'd150};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd174, 8'd164, 8'd163};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd154};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd168, 8'd159, 8'd156};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd4, 8'd3, 8'd4};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd174, 8'd180, 8'd180};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd162, 8'd168, 8'd164};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd45, 8'd45, 8'd43};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd153};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd39, 8'd36, 8'd35};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd162};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd170, 8'd159, 8'd155};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd6, 8'd4, 8'd5};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd165, 8'd154, 8'd153};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd173, 8'd164, 8'd162};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd113, 8'd117, 8'd124};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd86, 8'd82, 8'd81};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd0, 8'd0, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd174, 8'd165, 8'd164};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd155};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd155};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd174, 8'd166, 8'd163};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd90};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd171, 8'd162, 8'd158};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd155};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd164, 8'd155, 8'd153};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd233, 8'd238, 8'd255};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd146, 8'd136, 8'd135};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd90, 8'd85, 8'd86};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd155, 8'd148, 8'd146};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd164, 8'd155, 8'd153};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd0, 8'd0, 8'd2};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd169, 8'd157, 8'd157};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd124, 8'd120, 8'd116};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd168, 8'd159, 8'd155};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd39, 8'd37, 8'd36};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd171, 8'd164, 8'd163};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd155};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd159};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd103, 8'd96, 8'd94};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd164, 8'd155, 8'd153};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd175, 8'd164, 8'd163};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd201, 8'd213, 8'd245};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd243};
					endcase
				end
				`ybit'd12: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd238};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd235};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd188, 8'd201, 8'd223};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd174, 8'd190, 8'd200};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd162, 8'd177, 8'd179};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd153, 8'd170, 8'd169};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd148, 8'd166, 8'd158};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd142, 8'd160, 8'd151};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd140, 8'd155, 8'd147};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd143, 8'd157, 8'd151};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd145, 8'd158, 8'd152};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd146, 8'd157, 8'd153};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd150, 8'd160, 8'd154};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd155, 8'd170, 8'd165};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd167, 8'd181, 8'd182};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd202};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd183, 8'd197, 8'd213};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd205};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd161, 8'd177, 8'd176};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd148, 8'd164, 8'd153};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd142, 8'd160, 8'd147};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd143, 8'd160, 8'd148};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd147, 8'd163, 8'd155};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd153, 8'd169, 8'd166};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd157, 8'd171, 8'd171};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd157, 8'd172, 8'd171};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd154, 8'd168, 8'd167};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd149, 8'd165, 8'd155};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd146, 8'd161, 8'd149};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd145, 8'd159, 8'd147};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd150, 8'd164, 8'd155};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd159, 8'd171, 8'd171};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd169, 8'd182, 8'd189};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd183, 8'd195, 8'd211};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd189, 8'd200, 8'd224};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd191, 8'd203, 8'd227};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd192, 8'd204, 8'd227};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd216};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd170, 8'd183, 8'd192};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd159, 8'd171, 8'd172};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd155, 8'd164, 8'd163};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd153, 8'd163, 8'd159};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd153, 8'd164, 8'd155};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd149, 8'd162, 8'd149};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd146, 8'd159, 8'd142};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd144, 8'd156, 8'd144};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd143, 8'd156, 8'd144};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd149, 8'd153, 8'd147};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd64, 8'd56, 8'd59};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd127, 8'd119, 8'd117};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd143, 8'd135, 8'd132};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd42};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd10, 8'd10, 8'd9};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd65, 8'd62, 8'd61};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd152, 8'd143, 8'd142};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd174, 8'd164, 8'd163};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd153};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd171, 8'd160, 8'd159};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd159};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd155, 8'd145, 8'd143};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd2};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd153};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd159, 8'd149, 8'd147};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd82, 8'd79, 8'd77};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd88, 8'd85, 8'd83};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd79, 8'd72, 8'd72};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd190, 8'd180, 8'd179};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd172, 8'd162, 8'd159};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd154};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd31, 8'd28, 8'd28};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd27};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd27};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd21, 8'd18, 8'd17};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd89};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd167, 8'd158, 8'd155};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd152};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd129, 8'd121, 8'd119};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd31, 8'd28, 8'd27};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd28};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd33, 8'd31, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd219, 8'd223, 8'd235};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd156};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd144, 8'd134, 8'd133};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd174, 8'd164, 8'd163};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd54, 8'd47, 8'd47};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd95, 8'd89, 8'd89};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd88};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd168, 8'd156, 8'd155};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd32, 8'd28, 8'd28};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd174, 8'd166, 8'd164};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd57, 8'd52, 8'd50};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd98};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd1};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd175, 8'd165, 8'd163};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd28};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd17, 8'd17, 8'd16};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd32, 8'd29, 8'd28};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd15, 8'd14, 8'd14};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd27, 8'd26, 8'd25};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd28};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd169, 8'd163, 8'd160};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd155};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd173, 8'd164, 8'd162};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd32, 8'd29, 8'd28};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd28, 8'd24, 8'd24};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd200, 8'd213, 8'd243};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd242};
					endcase
				end
				`ybit'd13: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd195, 8'd206, 8'd234};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd233};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd191, 8'd203, 8'd225};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd180, 8'd195, 8'd212};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd172, 8'd186, 8'd199};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd165, 8'd179, 8'd187};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd158, 8'd173, 8'd176};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd150, 8'd163, 8'd161};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd146, 8'd157, 8'd154};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd149, 8'd157, 8'd158};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd153, 8'd160, 8'd162};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd150, 8'd157, 8'd160};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd150, 8'd158, 8'd160};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd157, 8'd168, 8'd168};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd168, 8'd178, 8'd185};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd174, 8'd187, 8'd197};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd178, 8'd189, 8'd201};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd171, 8'd184, 8'd193};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd156, 8'd171, 8'd167};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd145, 8'd161, 8'd150};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd140, 8'd156, 8'd145};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd142, 8'd154, 8'd145};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd143, 8'd155, 8'd146};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd145, 8'd160, 8'd151};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd148, 8'd163, 8'd157};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd150, 8'd165, 8'd159};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd148, 8'd163, 8'd157};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd145, 8'd161, 8'd149};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd141, 8'd155, 8'd142};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd139, 8'd151, 8'd141};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd143, 8'd156, 8'd146};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd148, 8'd161, 8'd153};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd159, 8'd173, 8'd174};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd170, 8'd183, 8'd191};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd205};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd179, 8'd193, 8'd206};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd182, 8'd195, 8'd212};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd178, 8'd190, 8'd205};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd168, 8'd181, 8'd188};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd164, 8'd170, 8'd173};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd159, 8'd164, 8'd165};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd156, 8'd162, 8'd161};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd155, 8'd161, 8'd154};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd153, 8'd159, 8'd151};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd149, 8'd157, 8'd147};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd147, 8'd154, 8'd143};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd148, 8'd155, 8'd144};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd82};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd167, 8'd159, 8'd153};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd39, 8'd37, 8'd36};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd173, 8'd164, 8'd164};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd159};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd168, 8'd157, 8'd155};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd169, 8'd158, 8'd156};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd175, 8'd167, 8'd165};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd39, 8'd38, 8'd36};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd164, 8'd157, 8'd152};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd172, 8'd161, 8'd159};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd88};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd178, 8'd165, 8'd165};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd1};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd163, 8'd153, 8'd151};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd157, 8'd147, 8'd146};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd169, 8'd161, 8'd158};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd1};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd88};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd163, 8'd154, 8'd153};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd166, 8'd159, 8'd156};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd88};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd128, 8'd128, 8'd128};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd80};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd97};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd153};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd172, 8'd166, 8'd164};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd88};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd149};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd141, 8'd133, 8'd132};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd27};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd112, 8'd107, 8'd107};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd153, 8'd148, 8'd145};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd161};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd158, 8'd156};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd2};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd94, 8'd90, 8'd89};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd170, 8'd159, 8'd154};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd7, 8'd3, 8'd6};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd199, 8'd206, 8'd230};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd238};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
					endcase
				end
				`ybit'd14: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd226};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd190, 8'd202, 8'd229};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd229};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd188, 8'd200, 8'd226};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd182, 8'd195, 8'd214};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd173, 8'd188, 8'd203};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd169, 8'd178, 8'd188};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd158, 8'd167, 8'd172};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd154, 8'd158, 8'd156};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd152, 8'd159, 8'd161};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd155, 8'd161, 8'd169};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd155, 8'd158, 8'd161};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd153, 8'd157, 8'd160};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd157, 8'd165, 8'd173};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd165, 8'd174, 8'd182};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd169, 8'd178, 8'd187};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd168, 8'd178, 8'd185};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd164, 8'd173, 8'd180};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd153, 8'd163, 8'd164};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd145, 8'd156, 8'd148};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd141, 8'd152, 8'd144};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd141, 8'd152, 8'd144};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd142, 8'd153, 8'd145};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd143, 8'd155, 8'd145};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd144, 8'd157, 8'd148};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd148, 8'd160, 8'd153};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd147, 8'd160, 8'd152};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd141, 8'd157, 8'd146};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd138, 8'd152, 8'd135};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd137, 8'd149, 8'd139};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd138, 8'd150, 8'd140};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd144, 8'd154, 8'd147};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd151, 8'd163, 8'd160};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd161, 8'd175, 8'd175};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd170, 8'd183, 8'd191};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd172, 8'd184, 8'd193};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd173, 8'd185, 8'd198};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd173, 8'd183, 8'd197};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd171, 8'd181, 8'd188};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd167, 8'd170, 8'd176};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd165, 8'd163, 8'd168};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd162, 8'd162, 8'd162};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd158, 8'd158, 8'd158};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd155, 8'd159, 8'd153};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd152, 8'd155, 8'd148};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd152, 8'd155, 8'd149};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd153, 8'd156, 8'd149};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd93, 8'd89, 8'd88};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd161};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd144, 8'd134, 8'd132};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd145, 8'd135, 8'd135};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd142, 8'd132, 8'd132};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd128, 8'd118, 8'd119};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd99, 8'd93, 8'd92};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd121, 8'd116, 8'd113};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd163, 8'd156, 8'd151};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd130, 8'd125, 8'd122};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd85};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd168, 8'd157, 8'd156};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd151};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd151, 8'd141, 8'd139};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd2};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd154};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd147, 8'd136, 8'd133};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd77};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd144, 8'd137, 8'd133};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd82, 8'd78, 8'd77};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd92, 8'd88, 8'd88};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd153};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd46, 8'd44, 8'd42};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd0};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd126, 8'd127, 8'd128};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd164, 8'd155, 8'd153};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd143, 8'd133, 8'd130};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd161, 8'd151, 8'd150};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd143, 8'd133, 8'd131};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd159};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd28, 8'd27, 8'd26};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd66};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd177, 8'd167, 8'd165};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd4};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd171, 8'd162, 8'd160};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd165, 8'd154, 8'd152};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd7, 8'd5, 8'd5};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd175, 8'd165, 8'd164};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd170, 8'd159, 8'd158};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd145, 8'd135, 8'd133};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd148, 8'd138, 8'd137};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd148, 8'd138, 8'd136};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd150, 8'd141, 8'd139};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd40};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd151};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd84};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd198, 8'd210, 8'd241};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd240};
					endcase
				end
				`ybit'd15: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd180, 8'd192, 8'd213};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd184, 8'd196, 8'd219};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd189, 8'd201, 8'd224};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd190, 8'd202, 8'd228};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd223};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd175, 8'd190, 8'd205};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd170, 8'd179, 8'd188};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd162, 8'd167, 8'd169};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd156, 8'd160, 8'd159};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd155, 8'd158, 8'd157};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd156, 8'd159, 8'd164};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd152, 8'd156, 8'd159};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd150, 8'd154, 8'd157};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd154, 8'd158, 8'd162};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd159, 8'd163, 8'd167};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd160, 8'd165, 8'd170};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd159, 8'd165, 8'd168};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd157, 8'd161, 8'd164};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd151, 8'd156, 8'd153};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd147, 8'd153, 8'd146};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd145, 8'd150, 8'd144};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd143, 8'd149, 8'd143};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd143, 8'd149, 8'd143};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd145, 8'd152, 8'd144};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd147, 8'd154, 8'd147};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd147, 8'd155, 8'd146};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd147, 8'd155, 8'd146};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd141, 8'd152, 8'd142};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd140, 8'd147, 8'd139};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd137, 8'd145, 8'd136};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd137, 8'd145, 8'd136};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd139, 8'd149, 8'd141};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd146, 8'd158, 8'd155};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd155, 8'd169, 8'd170};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd162, 8'd175, 8'd183};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd164, 8'd177, 8'd182};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd165, 8'd178, 8'd186};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd170, 8'd180, 8'd192};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd170, 8'd181, 8'd187};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd168, 8'd172, 8'd178};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd166, 8'd165, 8'd169};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd162, 8'd162, 8'd162};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd159, 8'd158, 8'd158};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd157, 8'd157, 8'd153};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd156, 8'd156, 8'd151};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd155, 8'd155, 8'd150};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd154, 8'd154, 8'd149};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd201, 8'd194, 8'd195};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd152};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd165, 8'd154, 8'd152};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd139};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd67, 8'd66, 8'd65};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd163, 8'd156, 8'd151};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd89, 8'd85, 8'd83};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd153, 8'd148, 8'd146};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd166, 8'd154, 8'd154};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd134};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd154};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd154};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd153};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd118, 8'd112, 8'd112};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd153};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd95, 8'd91, 8'd90};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd85, 8'd81, 8'd81};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd152};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd84};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd0};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd112, 8'd118, 8'd127};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd158, 8'd148, 8'd147};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd151, 8'd147, 8'd145};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd66, 8'd63, 8'd61};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd139, 8'd130, 8'd129};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd164};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd88};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd172, 8'd163, 8'd161};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd174, 8'd164, 8'd163};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd151};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd165, 8'd159, 8'd155};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd201, 8'd211, 8'd240};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd239};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd197, 8'd208, 8'd238};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd197, 8'd208, 8'd238};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
					endcase
				end
				`ybit'd16: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd172, 8'd184, 8'd198};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd177, 8'd192, 8'd208};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd182, 8'd197, 8'd220};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd185, 8'd200, 8'd222};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd181, 8'd195, 8'd213};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd173, 8'd185, 8'd195};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd165, 8'd174, 8'd174};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd159, 8'd166, 8'd162};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd154, 8'd159, 8'd154};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd151, 8'd156, 8'd154};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd150, 8'd155, 8'd154};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd151, 8'd152, 8'd154};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd148, 8'd149, 8'd150};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd149, 8'd150, 8'd154};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd151, 8'd152, 8'd156};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd149, 8'd153, 8'd152};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd149, 8'd153, 8'd153};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd150, 8'd152, 8'd149};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd149, 8'd150, 8'd147};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd149, 8'd151, 8'd146};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd149, 8'd150, 8'd146};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd147, 8'd148, 8'd143};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd145, 8'd148, 8'd142};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd144, 8'd149, 8'd142};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd146, 8'd151, 8'd144};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd146, 8'd152, 8'd144};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd145, 8'd151, 8'd143};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd140, 8'd149, 8'd140};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd137, 8'd145, 8'd138};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd136, 8'd142, 8'd137};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd136, 8'd141, 8'd137};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd137, 8'd144, 8'd140};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd144, 8'd151, 8'd147};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd152, 8'd162, 8'd162};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd159, 8'd169, 8'd175};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd161, 8'd172, 8'd174};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd163, 8'd174, 8'd177};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd167, 8'd177, 8'd186};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd169, 8'd178, 8'd188};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd168, 8'd171, 8'd177};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd164, 8'd165, 8'd169};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd160, 8'd160, 8'd160};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd157, 8'd157, 8'd157};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd155, 8'd154, 8'd150};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd158, 8'd155, 8'd150};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd159, 8'd155, 8'd152};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd169, 8'd164, 8'd161};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd156};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd162};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd157};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd179, 8'd170, 8'd168};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd159, 8'd151, 8'd145};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd182, 8'd177, 8'd173};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd169, 8'd158, 8'd156};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd84};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd130, 8'd120, 8'd119};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd157};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd5, 8'd4, 8'd4};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd177, 8'd167, 8'd164};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd155};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd170, 8'd162, 8'd158};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd153};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd165, 8'd158, 8'd152};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd170, 8'd165, 8'd161};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd121, 8'd116, 8'd113};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd171, 8'd165, 8'd162};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd40};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd85};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd159};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd96, 8'd98, 8'd104};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd172, 8'd178, 8'd199};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd174, 8'd180, 8'd207};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd175, 8'd181, 8'd205};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd144};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd159};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd172, 8'd166, 8'd164};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd170, 8'd159, 8'd158};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd157};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd156};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd153};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd121, 8'd119};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd90};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd154};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd169, 8'd162, 8'd160};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd54, 8'd50, 8'd51};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd171, 8'd165, 8'd162};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd174, 8'd167, 8'd164};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd171, 8'd162, 8'd160};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd246};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd197, 8'd207, 8'd237};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd237};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd195, 8'd206, 8'd236};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd231};
					endcase
				end
				`ybit'd17: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd166, 8'd179, 8'd188};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd169, 8'd185, 8'd196};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd174, 8'd190, 8'd207};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd175, 8'd191, 8'd207};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd171, 8'd186, 8'd200};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd164, 8'd178, 8'd184};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd158, 8'd167, 8'd160};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd158, 8'd160, 8'd153};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd154, 8'd155, 8'd148};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd151, 8'd152, 8'd147};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd149, 8'd149, 8'd144};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd143};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd141};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd147, 8'd144, 8'd145};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd145};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd144, 8'd144, 8'd144};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd144, 8'd144, 8'd141};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd142};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd143};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd145};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd151, 8'd148, 8'd145};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd142};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd141};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd145, 8'd147, 8'd140};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd146, 8'd147, 8'd141};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd148, 8'd148, 8'd143};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd145, 8'd147, 8'd140};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd143, 8'd146, 8'd139};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd140, 8'd143, 8'd137};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd136};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd138, 8'd138, 8'd136};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd138, 8'd140, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd143, 8'd146, 8'd144};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd150, 8'd156, 8'd157};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd156, 8'd161, 8'd169};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd157, 8'd168, 8'd170};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd158, 8'd169, 8'd172};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd163, 8'd174, 8'd179};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd163, 8'd174, 8'd179};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd163, 8'd167, 8'd172};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd159, 8'd160, 8'd164};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd158, 8'd158, 8'd157};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd155, 8'd155, 8'd154};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd154, 8'd153, 8'd149};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd156, 8'd153, 8'd148};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd158, 8'd154, 8'd151};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd85};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd173, 8'd162, 8'd161};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd155};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd89, 8'd85, 8'd85};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd89};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd85, 8'd82, 8'd80};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd132, 8'd127, 8'd124};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd168, 8'd157, 8'd155};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd6, 8'd6, 8'd5};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd173, 8'd164, 8'd163};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd157};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd159};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd0, 8'd0, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd141, 8'd134, 8'd134};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd102, 8'd95, 8'd95};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd147, 8'd137, 8'd136};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd2};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd154, 8'd144, 8'd142};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd159};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd175, 8'd167, 8'd164};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd169, 8'd160, 8'd155};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd153, 8'd146, 8'd145};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd3, 8'd0, 8'd1};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd4, 8'd0, 8'd1};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd0, 8'd0, 8'd1};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd89};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd167, 8'd158, 8'd156};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd105, 8'd108, 8'd115};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd185, 8'd201, 8'd219};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd189, 8'd204, 8'd230};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd191, 8'd205, 8'd235};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd208, 8'd217, 8'd243};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd163};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd144, 8'd134, 8'd133};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd142, 8'd132, 8'd131};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd139, 8'd129, 8'd128};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd169, 8'd164, 8'd162};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd153};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd175, 8'd168, 8'd166};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd68, 8'd65, 8'd64};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd94, 8'd93, 8'd90};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd1};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd107};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd0, 8'd2, 8'd1};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd170, 8'd167, 8'd162};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd181, 8'd176, 8'd173};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd149};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd111, 8'd114, 8'd124};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd190, 8'd208, 8'd232};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd187, 8'd199, 8'd222};
					endcase
				end
				`ybit'd18: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd160, 8'd173, 8'd179};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd160, 8'd176, 8'd183};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd162, 8'd180, 8'd186};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd162, 8'd180, 8'd187};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd158, 8'd175, 8'd179};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd154, 8'd166, 8'd166};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd152, 8'd159, 8'd154};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd154, 8'd157, 8'd150};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd153, 8'd154, 8'd146};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd149, 8'd150, 8'd144};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd147, 8'd147, 8'd141};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd147, 8'd143, 8'd140};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd145, 8'd141, 8'd140};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd139};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd139};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd139};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd139};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd138};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd140};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd149, 8'd146, 8'd141};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd152, 8'd149, 8'd144};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd149, 8'd146, 8'd141};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd139};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd145, 8'd144, 8'd139};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd146, 8'd145, 8'd140};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd145, 8'd146, 8'd140};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd145, 8'd146, 8'd140};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd144, 8'd145, 8'd140};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd138};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd135};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd135};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd137};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd140, 8'd141, 8'd141};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd144, 8'd148, 8'd150};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd150, 8'd154, 8'd157};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd150, 8'd159, 8'd160};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd153, 8'd161, 8'd163};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd155, 8'd166, 8'd168};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd155, 8'd165, 8'd167};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd152, 8'd161, 8'd160};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd152, 8'd158, 8'd156};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd153, 8'd154, 8'd152};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd151, 8'd151, 8'd149};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd152, 8'd151, 8'd147};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd154, 8'd151, 8'd146};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd156, 8'd153, 8'd146};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd87};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd163, 8'd155, 8'd153};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd64, 8'd57, 8'd55};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd17, 8'd17, 8'd17};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd174, 8'd168, 8'd169};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd168, 8'd161, 8'd155};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd3};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd177, 8'd168, 8'd166};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd2};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd169, 8'd159, 8'd157};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd154};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd4, 8'd3, 8'd3};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd164, 8'd155, 8'd153};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd163, 8'd160, 8'd158};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd2};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd147, 8'd139, 8'd137};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd156, 8'd151, 8'd148};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd176, 8'd166, 8'd165};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd38, 8'd37, 8'd35};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd162, 8'd155, 8'd150};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd156};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd100, 8'd95, 8'd93};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd25, 8'd23, 8'd23};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd25, 8'd23, 8'd22};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd25, 8'd23, 8'd22};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd15, 8'd14, 8'd14};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd89};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd66, 8'd59, 8'd60};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd43, 8'd44, 8'd48};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd44, 8'd45, 8'd50};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd45, 8'd45, 8'd51};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd132, 8'd138, 8'd144};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd165};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd142, 8'd132, 8'd131};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd89, 8'd78, 8'd82};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd170, 8'd159, 8'd157};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd154};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd1};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd153};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd146, 8'd136, 8'd138};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd110, 8'd99, 8'd102};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd125};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd3, 8'd2, 8'd3};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd163};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd0};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd196, 8'd202, 8'd225};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd120, 8'd125, 8'd142};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd80};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd165, 8'd158, 8'd155};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd42, 8'd40, 8'd39};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd236};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd235};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd182, 8'd193, 8'd215};
					endcase
				end
				`ybit'd19: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd152, 8'd166, 8'd167};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd148, 8'd166, 8'd165};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd147, 8'd166, 8'd164};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd146, 8'd165, 8'd162};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd144, 8'd163, 8'd158};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd143, 8'd157, 8'd150};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd147, 8'd154, 8'd146};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd149, 8'd151, 8'd145};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd149, 8'd150, 8'd143};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd147, 8'd148, 8'd142};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd144, 8'd144, 8'd138};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd137};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd144, 8'd139, 8'd138};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd138};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd138};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd136};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd137};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd142, 8'd140, 8'd136};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd137};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd147, 8'd144, 8'd139};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd148, 8'd145, 8'd140};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd147, 8'd144, 8'd139};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd136};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd137};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd145, 8'd144, 8'd139};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd143, 8'd144, 8'd138};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd143, 8'd144, 8'd138};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd142, 8'd142, 8'd138};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd138};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd136};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd135};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd137};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd141, 8'd138, 8'd139};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd142};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd147, 8'd147, 8'd147};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd148, 8'd150, 8'd149};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd147, 8'd156, 8'd155};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd148, 8'd159, 8'd156};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd147, 8'd159, 8'd155};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd145, 8'd154, 8'd149};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd147, 8'd153, 8'd147};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd149, 8'd150, 8'd144};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd148, 8'd149, 8'd143};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd149, 8'd148, 8'd143};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd153, 8'd150, 8'd145};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd154, 8'd151, 8'd146};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd168, 8'd163, 8'd161};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd148, 8'd139, 8'd137};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd126, 8'd118, 8'd115};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd18, 8'd14, 8'd15};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd31, 8'd27, 8'd31};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd17, 8'd15, 8'd18};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd154};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd153};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd155};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd0};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd174, 8'd163, 8'd161};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd154};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd160};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd153};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd154};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd175, 8'd167, 8'd163};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd37, 8'd34, 8'd34};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd168, 8'd155, 8'd152};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd155};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd134, 8'd126, 8'd124};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd92, 8'd88, 8'd87};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd167, 8'd157, 8'd153};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd169, 8'd160, 8'd158};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd166, 8'd156, 8'd152};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd168, 8'd155, 8'd153};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd150, 8'd138, 8'd135};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd163, 8'd153, 8'd151};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd93, 8'd89, 8'd89};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd88};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd167, 8'd158, 8'd156};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd164, 8'd154, 8'd152};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd164, 8'd156, 8'd152};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd160};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd155, 8'd148, 8'd146};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd155};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd119, 8'd121, 8'd127};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd175, 8'd165, 8'd163};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd172, 8'd162, 8'd161};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd152};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd1, 8'd2, 8'd1};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd158};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd153};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd167, 8'd159, 8'd156};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd2};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd155};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd168, 8'd158, 8'd156};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd167, 8'd156, 8'd154};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd2};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd167, 8'd158, 8'd154};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd165, 8'd156, 8'd153};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd165, 8'd157, 8'd155};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd165, 8'd155, 8'd153};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd158};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd169, 8'd160, 8'd156};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd1};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd3};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd190, 8'd205, 8'd231};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd207, 8'd216, 8'd240};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd18, 8'd17, 8'd18};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd5, 8'd3, 8'd3};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd166, 8'd155, 8'd151};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd167, 8'd158, 8'd154};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd131, 8'd123, 8'd120};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd235};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd235};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd232};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd190, 8'd202, 8'd231};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd188, 8'd200, 8'd229};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd188, 8'd201, 8'd229};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd188, 8'd200, 8'd230};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd189, 8'd199, 8'd229};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd228};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd187, 8'd199, 8'd228};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd189, 8'd201, 8'd230};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd231};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd231};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd189, 8'd200, 8'd230};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd231};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd228};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd179, 8'd192, 8'd212};
					endcase
				end
				`ybit'd20: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd144, 8'd160, 8'd154};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd138, 8'd158, 8'd148};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd134, 8'd154, 8'd143};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd132, 8'd152, 8'd142};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd132, 8'd152, 8'd141};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd134, 8'd150, 8'd140};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd140, 8'd149, 8'd141};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd146, 8'd148, 8'd142};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd147, 8'd148, 8'd142};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd146, 8'd145, 8'd141};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd137};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd138};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd142, 8'd137, 8'd134};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd134};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd136};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd136};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd136};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd145, 8'd142, 8'd137};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd138};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd145, 8'd142, 8'd137};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd135};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd135};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd138};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd137};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd139};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd137};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd135};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd135};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd140, 8'd138, 8'd139};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd142, 8'd140, 8'd141};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd143};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd145, 8'd145, 8'd143};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd144, 8'd148, 8'd143};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd144, 8'd150, 8'd145};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd143, 8'd149, 8'd145};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd143, 8'd150, 8'd143};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd144, 8'd149, 8'd143};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd146, 8'd147, 8'd142};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd145, 8'd146, 8'd141};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd146, 8'd145, 8'd140};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd151, 8'd148, 8'd143};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd163, 8'd158, 8'd154};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd171, 8'd165, 8'd160};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd172, 8'd161, 8'd158};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd161, 8'd156, 8'd153};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd2};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd10, 8'd8, 8'd11};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd24, 8'd20, 8'd22};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd157};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd174, 8'd163, 8'd159};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd154, 8'd150, 8'd149};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd11, 8'd10, 8'd10};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd168, 8'd162, 8'd158};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd79, 8'd76, 8'd74};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd167, 8'd163, 8'd159};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd43, 8'd41, 8'd40};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd171, 8'd164, 8'd159};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd158, 8'd150, 8'd146};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd133, 8'd128, 8'd129};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd88};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd156};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd94, 8'd91, 8'd91};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd94, 8'd91, 8'd89};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd88};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd159, 8'd154, 8'd151};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd83};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd169, 8'd162, 8'd156};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd167, 8'd161, 8'd158};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd85};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd167, 8'd161, 8'd156};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd86};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd88, 8'd85, 8'd84};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd175, 8'd164, 8'd163};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd36, 8'd33, 8'd31};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd165, 8'd157, 8'd152};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd170, 8'd162, 8'd158};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd75};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd157};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd111, 8'd114, 8'd118};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd108, 8'd102, 8'd101};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd169, 8'd161, 8'd161};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd175, 8'd164, 8'd160};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd172, 8'd166, 8'd161};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd141, 8'd135, 8'd130};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd170, 8'd162, 8'd157};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd0, 8'd0, 8'd0};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd176, 8'd165, 8'd162};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd172, 8'd162, 8'd158};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd169, 8'd163, 8'd160};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd175, 8'd164, 8'd161};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd174, 8'd163, 8'd160};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd171, 8'd160, 8'd159};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd0, 8'd1, 8'd2};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd174, 8'd164, 8'd160};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd172, 8'd161, 8'd158};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd172, 8'd161, 8'd160};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd183, 8'd188, 8'd208};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd184, 8'd187, 8'd219};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd231};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd192, 8'd201, 8'd236};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd171, 8'd165, 8'd162};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd170, 8'd160, 8'd156};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd172, 8'd164, 8'd158};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd205, 8'd214, 8'd240};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd232};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd189, 8'd201, 8'd228};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd226};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd187, 8'd199, 8'd226};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd222};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd185, 8'd195, 8'd221};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd183, 8'd193, 8'd217};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd183, 8'd193, 8'd216};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd181, 8'd191, 8'd214};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd183, 8'd189, 8'd214};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd181, 8'd191, 8'd214};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd181, 8'd191, 8'd215};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd184, 8'd194, 8'd218};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd222};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd221};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd221};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd184, 8'd196, 8'd221};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd184, 8'd196, 8'd221};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd224};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd227};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd193, 8'd204, 8'd234};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd192, 8'd203, 8'd233};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd181, 8'd193, 8'd217};
					endcase
				end
				`ybit'd21: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd138, 8'd151, 8'd146};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd130, 8'd152, 8'd137};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd128, 8'd149, 8'd135};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd126, 8'd147, 8'd133};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd128, 8'd146, 8'd134};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd130, 8'd146, 8'd135};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd136, 8'd145, 8'd137};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd142, 8'd146, 8'd139};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd145, 8'd145, 8'd141};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd146, 8'd142, 8'd139};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd142, 8'd138, 8'd135};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd133};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd140, 8'd135, 8'd132};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd139, 8'd135, 8'd132};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd139, 8'd135, 8'd132};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd133};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd134};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd142, 8'd138, 8'd135};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd142, 8'd140, 8'd135};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd141, 8'd139, 8'd136};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd136};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd137};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd138};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd139};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd138};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd136};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd135};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd135};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd140, 8'd138, 8'd139};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd138};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd139};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd140};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd141, 8'd144, 8'd140};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd138, 8'd143, 8'd139};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd139, 8'd144, 8'd140};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd143, 8'd146, 8'd140};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd144, 8'd145, 8'd140};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd144, 8'd144, 8'd139};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd137};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd144, 8'd143, 8'd139};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd149, 8'd145, 8'd141};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd156, 8'd148, 8'd148};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd30, 8'd27, 8'd26};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd31, 8'd28, 8'd31};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd0};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd8, 8'd6, 8'd8};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd31, 8'd29, 8'd31};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd1, 8'd1, 8'd1};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd44, 8'd43, 8'd45};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd3, 8'd2, 8'd2};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd15, 8'd14, 8'd16};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd2, 8'd0, 8'd1};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd83, 8'd83, 8'd82};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd28};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd17, 8'd19};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd18, 8'd16, 8'd18};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd3, 8'd2, 8'd3};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd28};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd17, 8'd15, 8'd17};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd28, 8'd26, 8'd28};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd17, 8'd16, 8'd18};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd17, 8'd16, 8'd17};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd29};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd17, 8'd15, 8'd18};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd20, 8'd18, 8'd21};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd31};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd108, 8'd112, 8'd108};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd31, 8'd28, 8'd31};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd20, 8'd17, 8'd21};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd30, 8'd27, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd16, 8'd15, 8'd17};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd26, 8'd24, 8'd27};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd1};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd29, 8'd26, 8'd29};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd32, 8'd30, 8'd32};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd2};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd31, 8'd29, 8'd31};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd231};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd230};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd230};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd187, 8'd199, 8'd228};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd5, 8'd3, 8'd5};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd17, 8'd16, 8'd17};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd33};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd28, 8'd27, 8'd24};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd189, 8'd202, 8'd231};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd190, 8'd200, 8'd233};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd189, 8'd200, 8'd230};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd189, 8'd200, 8'd230};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd228};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd186, 8'd200, 8'd226};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd224};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd184, 8'd198, 8'd223};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd183, 8'd196, 8'd221};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd183, 8'd193, 8'd217};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd179, 8'd190, 8'd213};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd176, 8'd187, 8'd208};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd175, 8'd183, 8'd204};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd175, 8'd181, 8'd200};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd173, 8'd179, 8'd198};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd170, 8'd179, 8'd196};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd171, 8'd178, 8'd193};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd170, 8'd178, 8'd193};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd173, 8'd180, 8'd196};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd176, 8'd184, 8'd204};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd177, 8'd188, 8'd211};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd177, 8'd188, 8'd209};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd173, 8'd184, 8'd205};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd174, 8'd185, 8'd205};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd175, 8'd186, 8'd206};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd179, 8'd190, 8'd210};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd184, 8'd194, 8'd219};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd188, 8'd197, 8'd227};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd190, 8'd200, 8'd233};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd189, 8'd200, 8'd230};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd190, 8'd201, 8'd231};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd184, 8'd195, 8'd223};
					endcase
				end
				`ybit'd22: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd134, 8'd148, 8'd138};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd127, 8'd148, 8'd133};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd125, 8'd146, 8'd131};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd125, 8'd146, 8'd131};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd127, 8'd145, 8'd133};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd128, 8'd145, 8'd134};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd135, 8'd145, 8'd136};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd140, 8'd144, 8'd137};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd144, 8'd143, 8'd139};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd137};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd138, 8'd134, 8'd131};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd137, 8'd133, 8'd130};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd129};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd129};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd138, 8'd134, 8'd131};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd132};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd133};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd133};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd134};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd134};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd136};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd141, 8'd139, 8'd135};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd136};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd137};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd139};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd138};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd135};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd135};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd135};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd135};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd141, 8'd137, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd139, 8'd137, 8'd138};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd138};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd138};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd138};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd141, 8'd141, 8'd139};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd139, 8'd139, 8'd137};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd140, 8'd140, 8'd137};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd140, 8'd142, 8'd137};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd141, 8'd142, 8'd136};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd136};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd145, 8'd141, 8'd138};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd153, 8'd143, 8'd144};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd149, 8'd146, 8'd145};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd25, 8'd23, 8'd24};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd0};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd1, 8'd0, 8'd2};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd125, 8'd120, 8'd116};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd23, 8'd22, 8'd23};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd5, 8'd3, 8'd4};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd16, 8'd15, 8'd17};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd15, 8'd13, 8'd14};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd29};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd2, 8'd1, 8'd1};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd174, 8'd174, 8'd163};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd31, 8'd29, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd31, 8'd29, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd3, 8'd1, 8'd2};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd29};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd22, 8'd21, 8'd23};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd25, 8'd23, 8'd26};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd5, 8'd3, 8'd6};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd16, 8'd15, 8'd17};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd31, 8'd29, 8'd32};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd61};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd166, 8'd170, 8'd162};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd30, 8'd27, 8'd31};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd100};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd28, 8'd26, 8'd29};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd5, 8'd3, 8'd4};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd38, 8'd36, 8'd39};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd11, 8'd9, 8'd12};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd17, 8'd16, 8'd16};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd14, 8'd13, 8'd15};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd16, 8'd14, 8'd15};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd27, 8'd25, 8'd28};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd100, 8'd105, 8'd115};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd182, 8'd194, 8'd216};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd180, 8'd193, 8'd214};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd181, 8'd193, 8'd214};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd181, 8'd193, 8'd215};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd13, 8'd14, 8'd16};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd18, 8'd19};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd17, 8'd15, 8'd16};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd180, 8'd185, 8'd207};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd184, 8'd195, 8'd225};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd186, 8'd197, 8'd225};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd228};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd223};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd185, 8'd198, 8'd223};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd183, 8'd196, 8'd221};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd183, 8'd195, 8'd217};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd185, 8'd194, 8'd216};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd184, 8'd192, 8'd213};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd179, 8'd189, 8'd205};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd177, 8'd187, 8'd202};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd175, 8'd183, 8'd197};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd172, 8'd179, 8'd193};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd169, 8'd176, 8'd188};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd167, 8'd172, 8'd183};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd165, 8'd172, 8'd181};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd163, 8'd170, 8'd178};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd163, 8'd168, 8'd177};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd163, 8'd166, 8'd177};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd164, 8'd167, 8'd178};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd167, 8'd169, 8'd181};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd168, 8'd173, 8'd188};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd169, 8'd176, 8'd190};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd167, 8'd174, 8'd186};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd165, 8'd173, 8'd184};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd165, 8'd173, 8'd183};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd167, 8'd174, 8'd186};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd172, 8'd179, 8'd195};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd180, 8'd186, 8'd208};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd184, 8'd194, 8'd219};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd186, 8'd197, 8'd226};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd228};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd228};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd185, 8'd196, 8'd226};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd224};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd186, 8'd198, 8'd223};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd223};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd228};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd229};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd226};
					endcase
				end
				`ybit'd23: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd133, 8'd142, 8'd133};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd127, 8'd144, 8'd133};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd125, 8'd144, 8'd132};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd125, 8'd144, 8'd130};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd128, 8'd144, 8'd133};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd128, 8'd144, 8'd133};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd133, 8'd142, 8'd134};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd138, 8'd143, 8'd136};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd142, 8'd142, 8'd136};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd130};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd133, 8'd133, 8'd128};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd133, 8'd134, 8'd129};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd129};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd130};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd130};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd138, 8'd134, 8'd131};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd131};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd129};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd134, 8'd134, 8'd129};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd136, 8'd136, 8'd130};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd131};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd131};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd142, 8'd138, 8'd135};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd139};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd145, 8'd139, 8'd141};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd140};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd137, 8'd135, 8'd137};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd141, 8'd133, 8'd134};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd138, 8'd134, 8'd133};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd137, 8'd133, 8'd132};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd135};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd134};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd134};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd134};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd134};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd136, 8'd137, 8'd132};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd137, 8'd138, 8'd133};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd136, 8'd137, 8'd132};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd139, 8'd140, 8'd135};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd139, 8'd140, 8'd134};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd133};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd133};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd132};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd145, 8'd138, 8'd136};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd141};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd152, 8'd148, 8'd146};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd80};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd34, 8'd32, 8'd33};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd4, 8'd2, 8'd3};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd72, 8'd69, 8'd67};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd146, 8'd137, 8'd132};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd141, 8'd132, 8'd126};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd25, 8'd27, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd29, 8'd29, 8'd32};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd5, 8'd4, 8'd6};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd2, 8'd2, 8'd4};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd29, 8'd29, 8'd31};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd29};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd4, 8'd2, 8'd3};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd29};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd17, 8'd16, 8'd18};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd159, 8'd159, 8'd149};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd14, 8'd13, 8'd15};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd51, 8'd49, 8'd52};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd28, 8'd28, 8'd31};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd12, 8'd10, 8'd10};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd29, 8'd29, 8'd33};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd31, 8'd27, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd31};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd31};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd33};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd17, 8'd17, 8'd17};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd65, 8'd66, 8'd59};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd9, 8'd8, 8'd8};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd29, 8'd28, 8'd27};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd30, 8'd29, 8'd28};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd31, 8'd30, 8'd29};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd29};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd28};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd153, 8'd159, 8'd140};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd17, 8'd15, 8'd16};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd15, 8'd13, 8'd14};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd9, 8'd8, 8'd9};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd79};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd31, 8'd28, 8'd27};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd31, 8'd27, 8'd27};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd14, 8'd12, 8'd14};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd17, 8'd15, 8'd20};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd31, 8'd27, 8'd31};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd107};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd60};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd87, 8'd89, 8'd91};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd30, 8'd27, 8'd31};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd37, 8'd34, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd31, 8'd28, 8'd32};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd169, 8'd183, 8'd196};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd167, 8'd182, 8'd193};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd166, 8'd180, 8'd190};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd166, 8'd180, 8'd190};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd169, 8'd178, 8'd192};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd96, 8'd102, 8'd106};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd15, 8'd13, 8'd16};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd31};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd90, 8'd93, 8'd97};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd168, 8'd181, 8'd199};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd172, 8'd185, 8'd210};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd177, 8'd190, 8'd215};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd214};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd176, 8'd188, 8'd211};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd174, 8'd187, 8'd204};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd172, 8'd186, 8'd199};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd175, 8'd187, 8'd199};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd178, 8'd187, 8'd199};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd175, 8'd184, 8'd196};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd170, 8'd178, 8'd189};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd168, 8'd176, 8'd183};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd164, 8'd172, 8'd179};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd162, 8'd169, 8'd176};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd161, 8'd166, 8'd171};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd159, 8'd164, 8'd169};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd158, 8'd163, 8'd167};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd156, 8'd161, 8'd165};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd156, 8'd161, 8'd167};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd155, 8'd158, 8'd164};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd158, 8'd161, 8'd167};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd159, 8'd162, 8'd168};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd159, 8'd161, 8'd171};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd156, 8'd162, 8'd170};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd155, 8'd160, 8'd169};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd156, 8'd160, 8'd169};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd158, 8'd161, 8'd170};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd160, 8'd162, 8'd172};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd165, 8'd169, 8'd179};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd170, 8'd179, 8'd193};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd175, 8'd186, 8'd207};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd215};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd180, 8'd193, 8'd218};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd182, 8'd194, 8'd220};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd182, 8'd193, 8'd222};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd178, 8'd190, 8'd217};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd177, 8'd189, 8'd210};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd177, 8'd189, 8'd210};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd178, 8'd191, 8'd212};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd180, 8'd193, 8'd216};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd180, 8'd193, 8'd218};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd180, 8'd192, 8'd218};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd180, 8'd192, 8'd218};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd182, 8'd193, 8'd222};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd184, 8'd195, 8'd224};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd184, 8'd195, 8'd224};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd185, 8'd197, 8'd224};
					endcase
				end
				`ybit'd24: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd136, 8'd139, 8'd132};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd129, 8'd141, 8'd131};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd129, 8'd141, 8'd131};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd131, 8'd143, 8'd132};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd127, 8'd145, 8'd127};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd129, 8'd146, 8'd129};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd133, 8'd143, 8'd128};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd137, 8'd142, 8'd128};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd140, 8'd140, 8'd134};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd131};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd128};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd128};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd132, 8'd133, 8'd128};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd129};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd129};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd129};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd129};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd129};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd128};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd129, 8'd133, 8'd127};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd129, 8'd136, 8'd122};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd132, 8'd136, 8'd128};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd133, 8'd137, 8'd129};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd137, 8'd138, 8'd133};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd140, 8'd141, 8'd138};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd140, 8'd141, 8'd140};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd138, 8'd138, 8'd139};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd137};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd133};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd133};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd133};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd133};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd132};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd133, 8'd135, 8'd132};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd133, 8'd135, 8'd132};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd133, 8'd136, 8'd132};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd134, 8'd135, 8'd130};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd136, 8'd137, 8'd132};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd136, 8'd137, 8'd132};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd136, 8'd137, 8'd132};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd136, 8'd137, 8'd131};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd133, 8'd136, 8'd126};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd133, 8'd136, 8'd125};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd134, 8'd134, 8'd125};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd132};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd138};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd149, 8'd145, 8'd144};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd152, 8'd148, 8'd147};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd22, 8'd21, 8'd23};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd24, 8'd22, 8'd24};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd25, 8'd23, 8'd24};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd136};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd146, 8'd136, 8'd132};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd140, 8'd133, 8'd126};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd135, 8'd127, 8'd121};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd27, 8'd22, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd25, 8'd20, 8'd19};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd21, 8'd18, 8'd17};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd73, 8'd69, 8'd67};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd23, 8'd23, 8'd21};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd23, 8'd22, 8'd22};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd137};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd23, 8'd21, 8'd22};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd30, 8'd29, 8'd28};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd36, 8'd35, 8'd34};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd160, 8'd160, 8'd150};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd92};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd25, 8'd24, 8'd23};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd27, 8'd23, 8'd22};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd89, 8'd82, 8'd79};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd21, 8'd19, 8'd18};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd26, 8'd21, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd25, 8'd20, 8'd19};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd25, 8'd20, 8'd20};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd26, 8'd20, 8'd19};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd25, 8'd22, 8'd20};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd22, 8'd18, 8'd17};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd84, 8'd84, 8'd72};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd23, 8'd22, 8'd19};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd24, 8'd23, 8'd20};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd21, 8'd21, 8'd17};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd23, 8'd22, 8'd21};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd23, 8'd23, 8'd21};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd22, 8'd22, 8'd20};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd143, 8'd150, 8'd126};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd23, 8'd25, 8'd23};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd21, 8'd23, 8'd22};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd22, 8'd17};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd77};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd23, 8'd24, 8'd21};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd23, 8'd25, 8'd22};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd81};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd21, 8'd18};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd23, 8'd24, 8'd28};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd24, 8'd25, 8'd29};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd159, 8'd172, 8'd188};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd23, 8'd24, 8'd29};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd23, 8'd24, 8'd26};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd21, 8'd22};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd98};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd23, 8'd25, 8'd23};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd23, 8'd25, 8'd22};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd83};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd151, 8'd164, 8'd165};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd153, 8'd165, 8'd156};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd153, 8'd165, 8'd156};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd153, 8'd165, 8'd156};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd152, 8'd165, 8'd156};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd163, 8'd173, 8'd166};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd23, 8'd26, 8'd23};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd24, 8'd26, 8'd23};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd80, 8'd83, 8'd80};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd148, 8'd160, 8'd154};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd155, 8'd165, 8'd168};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd159, 8'd168, 8'd178};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd162, 8'd171, 8'd184};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd164, 8'd174, 8'd183};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd165, 8'd173, 8'd185};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd162, 8'd172, 8'd176};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd159, 8'd170, 8'd169};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd163, 8'd172, 8'd172};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd169, 8'd175, 8'd175};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd167, 8'd172, 8'd172};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd163, 8'd167, 8'd165};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd160, 8'd164, 8'd163};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd156, 8'd160, 8'd160};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd155, 8'd159, 8'd159};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd154, 8'd159, 8'd161};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd152, 8'd158, 8'd159};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd153, 8'd159, 8'd156};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd152, 8'd158, 8'd156};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd150, 8'd156, 8'd157};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd151, 8'd155, 8'd157};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd151, 8'd155, 8'd157};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd151, 8'd155, 8'd157};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd150, 8'd154, 8'd153};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd149, 8'd151, 8'd151};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd146, 8'd152, 8'd151};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd147, 8'd153, 8'd151};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd147, 8'd151, 8'd151};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd150, 8'd155, 8'd154};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd155, 8'd161, 8'd159};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd158, 8'd169, 8'd172};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd166, 8'd173, 8'd184};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd168, 8'd177, 8'd191};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd172, 8'd179, 8'd197};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd175, 8'd183, 8'd201};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd172, 8'd185, 8'd203};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd171, 8'd179, 8'd193};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd166, 8'd175, 8'd182};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd166, 8'd175, 8'd182};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd169, 8'd178, 8'd185};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd170, 8'd179, 8'd188};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd171, 8'd179, 8'd192};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd171, 8'd179, 8'd193};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd172, 8'd179, 8'd197};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd175, 8'd182, 8'd203};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd174, 8'd186, 8'd205};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd175, 8'd188, 8'd207};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd177, 8'd190, 8'd211};
					endcase
				end
				`ybit'd25: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd134, 8'd137, 8'd130};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd130, 8'd139, 8'd130};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd129, 8'd139, 8'd130};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd128, 8'd140, 8'd128};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd127, 8'd143, 8'd130};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd127, 8'd145, 8'd127};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd130, 8'd141, 8'd125};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd132, 8'd139, 8'd127};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd132, 8'd137, 8'd126};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd132, 8'd135, 8'd124};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd129, 8'd131, 8'd122};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd130, 8'd131, 8'd124};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd127, 8'd132, 8'd124};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd131, 8'd133, 8'd127};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd131, 8'd133, 8'd127};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd127};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd127};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd127};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd131, 8'd132, 8'd122};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd127, 8'd135, 8'd122};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd124, 8'd135, 8'd118};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd119};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd121};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd132, 8'd137, 8'd132};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd137, 8'd138, 8'd137};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd137, 8'd139, 8'd138};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd135, 8'd137, 8'd135};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd134, 8'd135, 8'd130};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd129};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd136, 8'd131, 8'd129};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd137, 8'd133, 8'd130};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd133, 8'd133, 8'd128};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd131, 8'd132, 8'd126};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd129, 8'd131, 8'd123};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd128, 8'd130, 8'd123};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd123};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd129, 8'd132, 8'd125};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd126};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd132, 8'd133, 8'd128};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd133, 8'd135, 8'd126};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd130, 8'd136, 8'd121};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd127, 8'd133, 8'd119};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd127, 8'd132, 8'd118};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd129, 8'd132, 8'd121};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd132, 8'd132, 8'd126};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd134};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd144, 8'd143, 8'd139};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd147, 8'd146, 8'd144};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd147};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd149, 8'd146, 8'd145};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd148, 8'd144, 8'd143};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd138};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd142, 8'd137, 8'd132};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd139, 8'd130, 8'd125};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd136, 8'd127, 8'd122};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd136, 8'd127, 8'd122};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd137, 8'd128, 8'd123};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd138, 8'd128, 8'd126};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd138, 8'd129, 8'd126};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd136, 8'd131, 8'd127};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd135, 8'd131, 8'd129};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd135, 8'd133, 8'd134};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd135, 8'd133, 8'd133};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd138, 8'd138, 8'd136};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd149, 8'd149, 8'd142};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd163, 8'd161, 8'd149};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd166, 8'd163, 8'd150};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd158, 8'd154, 8'd142};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd148, 8'd139, 8'd129};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd142, 8'd132, 8'd121};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd141, 8'd131, 8'd119};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd143, 8'd131, 8'd119};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd141, 8'd129, 8'd117};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd140, 8'd128, 8'd114};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd141, 8'd129, 8'd115};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd139, 8'd131, 8'd116};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd138, 8'd131, 8'd115};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd130, 8'd133, 8'd111};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd111};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd111};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd111};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd111};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd130, 8'd132, 8'd110};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd110};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd127, 8'd135, 8'd111};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd129, 8'd139, 8'd112};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd131, 8'd141, 8'd114};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd131, 8'd141, 8'd114};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd130, 8'd140, 8'd113};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd130, 8'd141, 8'd116};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd135, 8'd142, 8'd124};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd139, 8'd147, 8'd143};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd139, 8'd151, 8'd159};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd138, 8'd150, 8'd159};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd138, 8'd151, 8'd152};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd136, 8'd149, 8'd139};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd136, 8'd149, 8'd139};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd138, 8'd148, 8'd137};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd136, 8'd147, 8'd132};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd137, 8'd148, 8'd132};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd138, 8'd150, 8'd133};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd138, 8'd151, 8'd134};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd137, 8'd150, 8'd131};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd138, 8'd152, 8'd131};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd137, 8'd151, 8'd130};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd138, 8'd148, 8'd131};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd137, 8'd150, 8'd132};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd137, 8'd150, 8'd132};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd135, 8'd147, 8'd129};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd135, 8'd145, 8'd128};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd138, 8'd147, 8'd132};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd140, 8'd148, 8'd141};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd143, 8'd149, 8'd150};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd145, 8'd151, 8'd155};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd148, 8'd156, 8'd154};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd148, 8'd156, 8'd153};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd145, 8'd155, 8'd145};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd143, 8'd152, 8'd141};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd148, 8'd157, 8'd146};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd153, 8'd160, 8'd150};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd153, 8'd159, 8'd149};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd153, 8'd155, 8'd146};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd149, 8'd152, 8'd145};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd147, 8'd152, 8'd144};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd146, 8'd151, 8'd149};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd146, 8'd154, 8'd147};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd147, 8'd154, 8'd148};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd147, 8'd154, 8'd147};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd146, 8'd154, 8'd146};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd145, 8'd152, 8'd145};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd146, 8'd151, 8'd145};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd146, 8'd151, 8'd145};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd145, 8'd150, 8'd144};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd141, 8'd147, 8'd140};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd141, 8'd146, 8'd139};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd141, 8'd146, 8'd137};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd141, 8'd146, 8'd138};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd141, 8'd146, 8'd138};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd141, 8'd147, 8'd140};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd145, 8'd152, 8'd144};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd149, 8'd156, 8'd148};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd151, 8'd159, 8'd157};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd153, 8'd161, 8'd161};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd157, 8'd164, 8'd170};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd162, 8'd169, 8'd174};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd160, 8'd169, 8'd176};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd156, 8'd167, 8'd166};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd152, 8'd163, 8'd157};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd151, 8'd162, 8'd156};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd152, 8'd164, 8'd158};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd153, 8'd165, 8'd161};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd154, 8'd164, 8'd165};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd152, 8'd163, 8'd164};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd156, 8'd166, 8'd169};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd159, 8'd168, 8'd174};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd161, 8'd171, 8'd177};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd165, 8'd174, 8'd181};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd167, 8'd175, 8'd187};
					endcase
				end
				`ybit'd26: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd130, 8'd132, 8'd126};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd131, 8'd134, 8'd128};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd130, 8'd135, 8'd128};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd131, 8'd139, 8'd128};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd128, 8'd138, 8'd126};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd125, 8'd140, 8'd122};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd127, 8'd138, 8'd122};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd124, 8'd137, 8'd119};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd123, 8'd135, 8'd118};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd124, 8'd134, 8'd116};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd113};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd115};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd118};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd121};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd127, 8'd135, 8'd123};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd126};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd126};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd126};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd120};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd117};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd122, 8'd134, 8'd116};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd119, 8'd132, 8'd114};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd121, 8'd134, 8'd117};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd124, 8'd134, 8'd122};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd128};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd133, 8'd137, 8'd130};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd132, 8'd135, 8'd128};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd132, 8'd133, 8'd125};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd132, 8'd133, 8'd124};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd131, 8'd132, 8'd124};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd131, 8'd132, 8'd123};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd128, 8'd133, 8'd122};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd127, 8'd129, 8'd116};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd120, 8'd128, 8'd112};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd118, 8'd126, 8'd111};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd119, 8'd125, 8'd111};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd115};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd119};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd120};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd119};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd123, 8'd136, 8'd114};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd120, 8'd132, 8'd111};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd119, 8'd131, 8'd110};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd114};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd124, 8'd131, 8'd117};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd133, 8'd133, 8'd127};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd135};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd143, 8'd141, 8'd139};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd143};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd142};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd146, 8'd142, 8'd140};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd144, 8'd140, 8'd137};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd141, 8'd136, 8'd134};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd126};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd132, 8'd128, 8'd121};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd135, 8'd126, 8'd121};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd134, 8'd125, 8'd120};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd135, 8'd125, 8'd123};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd135, 8'd126, 8'd123};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd133, 8'd128, 8'd124};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd127};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd132, 8'd130, 8'd131};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd133, 8'd131, 8'd132};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd134, 8'd134, 8'd132};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd145, 8'd145, 8'd138};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd159, 8'd158, 8'd145};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd163, 8'd161, 8'd148};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd157, 8'd153, 8'd141};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd135};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd142, 8'd131, 8'd126};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd141, 8'd130, 8'd124};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd142, 8'd130, 8'd118};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd139, 8'd127, 8'd115};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd139, 8'd128, 8'd114};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd140, 8'd127, 8'd114};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd141, 8'd127, 8'd114};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd136, 8'd128, 8'd113};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd135, 8'd128, 8'd113};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd134, 8'd128, 8'd113};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd133, 8'd129, 8'd114};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd135, 8'd128, 8'd114};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd134, 8'd128, 8'd110};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd132, 8'd127, 8'd109};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd132, 8'd125, 8'd111};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd130, 8'd126, 8'd108};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd127, 8'd130, 8'd108};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd127, 8'd131, 8'd108};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd130, 8'd135, 8'd110};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd130, 8'd136, 8'd110};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd129, 8'd134, 8'd109};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd128, 8'd133, 8'd108};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd127, 8'd132, 8'd109};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd131, 8'd133, 8'd114};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd135, 8'd139, 8'd127};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd133, 8'd142, 8'd140};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd129, 8'd144, 8'd138};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd131, 8'd141, 8'd132};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd130, 8'd144, 8'd122};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd129, 8'd144, 8'd121};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd130, 8'd142, 8'd118};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd130, 8'd142, 8'd113};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd129, 8'd142, 8'd114};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd130, 8'd142, 8'd115};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd130, 8'd140, 8'd114};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd130, 8'd140, 8'd113};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd129, 8'd140, 8'd111};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd130, 8'd141, 8'd111};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd132, 8'd139, 8'd113};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd131, 8'd141, 8'd114};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd130, 8'd140, 8'd113};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd139, 8'd112};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd130, 8'd138, 8'd111};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd130, 8'd135, 8'd112};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd130, 8'd134, 8'd118};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd130, 8'd133, 8'd124};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd132, 8'd135, 8'd124};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd135, 8'd139, 8'd125};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd135, 8'd141, 8'd124};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd134, 8'd140, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd134, 8'd140, 8'd119};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd137, 8'd142, 8'd122};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd142, 8'd145, 8'd126};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd142, 8'd145, 8'd126};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd124};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd128};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd142, 8'd143, 8'd127};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd143, 8'd144, 8'd133};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd142, 8'd145, 8'd136};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd140, 8'd148, 8'd137};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd140, 8'd149, 8'd135};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd140, 8'd149, 8'd134};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd140, 8'd148, 8'd130};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd140, 8'd147, 8'd133};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd140, 8'd147, 8'd133};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd137, 8'd144, 8'd129};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd136, 8'd143, 8'd125};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd123};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd133, 8'd139, 8'd124};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd133, 8'd139, 8'd124};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd133, 8'd139, 8'd125};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd134, 8'd142, 8'd124};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd135, 8'd144, 8'd125};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd140, 8'd148, 8'd130};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd141, 8'd146, 8'd132};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd141, 8'd146, 8'd133};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd144, 8'd148, 8'd141};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd148, 8'd152, 8'd146};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd149, 8'd156, 8'd147};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd155, 8'd141};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd143, 8'd152, 8'd135};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd142, 8'd151, 8'd133};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd141, 8'd150, 8'd133};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd140, 8'd149, 8'd133};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd139, 8'd147, 8'd135};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd140, 8'd148, 8'd136};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd142, 8'd150, 8'd139};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd146, 8'd152, 8'd144};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd148, 8'd155, 8'd147};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd152, 8'd158, 8'd150};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd155, 8'd161, 8'd154};
					endcase
				end
				`ybit'd27: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd126, 8'd129, 8'd122};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd127, 8'd131, 8'd122};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd122};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd121};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd124, 8'd135, 8'd119};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd117};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd121, 8'd133, 8'd116};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd118, 8'd133, 8'd112};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd117, 8'd132, 8'd111};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd117, 8'd129, 8'd109};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd116, 8'd128, 8'd109};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd117, 8'd128, 8'd111};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd119, 8'd131, 8'd114};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd118};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd119};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd125, 8'd132, 8'd121};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd126, 8'd129, 8'd123};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd127, 8'd130, 8'd123};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd118};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd113};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd117, 8'd132, 8'd111};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd115, 8'd130, 8'd109};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd115, 8'd129, 8'd113};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd120, 8'd131, 8'd117};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd125};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd131, 8'd134, 8'd127};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd129, 8'd132, 8'd125};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd120};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd118};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd126, 8'd131, 8'd118};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd118};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd123, 8'd129, 8'd116};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd120, 8'd128, 8'd111};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd116, 8'd125, 8'd105};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd114, 8'd123, 8'd103};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd114, 8'd123, 8'd103};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd116, 8'd125, 8'd106};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd119, 8'd125, 8'd111};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd121, 8'd128, 8'd114};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd115};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd120, 8'd132, 8'd110};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd118, 8'd130, 8'd106};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd116, 8'd127, 8'd104};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd117, 8'd126, 8'd106};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd123, 8'd127, 8'd109};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd128, 8'd130, 8'd116};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd133, 8'd134, 8'd126};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd138, 8'd139, 8'd133};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd139};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd139};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd138};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd140, 8'd136, 8'd133};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd135, 8'd130, 8'd126};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd132, 8'd127, 8'd123};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd133, 8'd124, 8'd119};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd133, 8'd124, 8'd119};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd131, 8'd125, 8'd119};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd130, 8'd125, 8'd120};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd132, 8'd127, 8'd123};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd133, 8'd130, 8'd124};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd129};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd129, 8'd126, 8'd128};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd130, 8'd131, 8'd125};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd138, 8'd140, 8'd127};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd148, 8'd149, 8'd133};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd152, 8'd153, 8'd137};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd136};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd130};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd139, 8'd131, 8'd126};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd139, 8'd131, 8'd125};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd140, 8'd130, 8'd120};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd140, 8'd128, 8'd116};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd139, 8'd125, 8'd112};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd139, 8'd125, 8'd112};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd139, 8'd125, 8'd112};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd137, 8'd125, 8'd113};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd133, 8'd124, 8'd112};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd134, 8'd126, 8'd113};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd134, 8'd125, 8'd113};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd133, 8'd125, 8'd112};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd130, 8'd122, 8'd109};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd130, 8'd122, 8'd109};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd130, 8'd122, 8'd109};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd127, 8'd124, 8'd107};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd125, 8'd127, 8'd106};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd127, 8'd129, 8'd108};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd129, 8'd130, 8'd110};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd129, 8'd130, 8'd107};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd107};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd105};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd126, 8'd128, 8'd110};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd129, 8'd134, 8'd117};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd127, 8'd138, 8'd119};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd127, 8'd139, 8'd120};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd128, 8'd140, 8'd117};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd127, 8'd140, 8'd111};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd127, 8'd140, 8'd111};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd125, 8'd138, 8'd109};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd126, 8'd136, 8'd109};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd108};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd127, 8'd136, 8'd109};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd108};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd128, 8'd133, 8'd110};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd108};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd125, 8'd135, 8'd108};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd108};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd127, 8'd136, 8'd109};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd110};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd109};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd126, 8'd131, 8'd108};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd126, 8'd129, 8'd108};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd107};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd123, 8'd125, 8'd111};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd122, 8'd125, 8'd109};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd110};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd110};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd109};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd128, 8'd130, 8'd109};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd112};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd133, 8'd131, 8'd112};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd133, 8'd131, 8'd112};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd116};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd136, 8'd134, 8'd118};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd136, 8'd133, 8'd124};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd133, 8'd136, 8'd124};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd132, 8'd138, 8'd123};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd131, 8'd139, 8'd123};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd133, 8'd141, 8'd124};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd123};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd123};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd123};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd132, 8'd139, 8'd121};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd131, 8'd139, 8'd118};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd130, 8'd138, 8'd117};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd117};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd126, 8'd133, 8'd115};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd127, 8'd134, 8'd116};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd127, 8'd136, 8'd115};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd130, 8'd138, 8'd116};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd118};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd134, 8'd139, 8'd122};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd133, 8'd135, 8'd122};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd133, 8'd137, 8'd122};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd136, 8'd141, 8'd125};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd138, 8'd145, 8'd128};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd137, 8'd147, 8'd123};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd137, 8'd147, 8'd123};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd134, 8'd144, 8'd121};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd133, 8'd142, 8'd122};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd138, 8'd120};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd120};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd120};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd131, 8'd138, 8'd122};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd125};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd137, 8'd143, 8'd127};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd141, 8'd148, 8'd130};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd144, 8'd150, 8'd135};
					endcase
				end
				`ybit'd28: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd120, 8'd123, 8'd115};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd123, 8'd127, 8'd117};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd122, 8'd129, 8'd115};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd120, 8'd132, 8'd115};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd114};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd118, 8'd128, 8'd112};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd116, 8'd127, 8'd110};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd114, 8'd127, 8'd108};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd113, 8'd128, 8'd107};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd111, 8'd128, 8'd106};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd112, 8'd130, 8'd108};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd113, 8'd130, 8'd106};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd115, 8'd130, 8'd107};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd116, 8'd131, 8'd112};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd117, 8'd132, 8'd112};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd119, 8'd129, 8'd114};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd122, 8'd129, 8'd119};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd123, 8'd129, 8'd120};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd116};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd120, 8'd132, 8'd112};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd115, 8'd130, 8'd108};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd113, 8'd126, 8'd106};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd113, 8'd126, 8'd108};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd117, 8'd126, 8'd113};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd119};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd126, 8'd129, 8'd122};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd126, 8'd129, 8'd122};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd116};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd123, 8'd130, 8'd113};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd115};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd120, 8'd128, 8'd112};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd120, 8'd128, 8'd109};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd103};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd112, 8'd124, 8'd98};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd97};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd111, 8'd121, 8'd98};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd111, 8'd121, 8'd100};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd103};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd115, 8'd125, 8'd106};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd117, 8'd128, 8'd106};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd116, 8'd128, 8'd106};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd116, 8'd127, 8'd103};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd113, 8'd124, 8'd100};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd114, 8'd124, 8'd99};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd117, 8'd125, 8'd102};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd121, 8'd127, 8'd108};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd125, 8'd130, 8'd116};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd131, 8'd136, 8'd123};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd136, 8'd138, 8'd130};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd139, 8'd141, 8'd136};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd139, 8'd140, 8'd135};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd139, 8'd137, 8'd134};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd129};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd137, 8'd129, 8'd125};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd133, 8'd125, 8'd120};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd130, 8'd124, 8'd116};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd130, 8'd123, 8'd116};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd129, 8'd123, 8'd116};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd130, 8'd124, 8'd118};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd133, 8'd126, 8'd121};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd133, 8'd128, 8'd124};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd128};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd126, 8'd126, 8'd126};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd128, 8'd129, 8'd121};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd133, 8'd135, 8'd119};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd138, 8'd138, 8'd122};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd124};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd141, 8'd138, 8'd128};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd136, 8'd133, 8'd126};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd123};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd136, 8'd131, 8'd124};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd139, 8'd130, 8'd120};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd139, 8'd126, 8'd115};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd136, 8'd124, 8'd112};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd135, 8'd123, 8'd111};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd135, 8'd122, 8'd110};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd135, 8'd123, 8'd110};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd135, 8'd123, 8'd111};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd135, 8'd123, 8'd111};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd134, 8'd122, 8'd110};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd130, 8'd121, 8'd109};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd129, 8'd121, 8'd108};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd129, 8'd121, 8'd108};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd127, 8'd119, 8'd106};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd126, 8'd121, 8'd105};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd122, 8'd124, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd125, 8'd126, 8'd108};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd131, 8'd126, 8'd109};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd130, 8'd125, 8'd108};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd128, 8'd122, 8'd108};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd127, 8'd121, 8'd106};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd127, 8'd121, 8'd106};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd106};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd105};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd108};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd123, 8'd136, 8'd107};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd123, 8'd138, 8'd109};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd124, 8'd136, 8'd105};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd124, 8'd136, 8'd106};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd122, 8'd136, 8'd104};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd105};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd104};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd105};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd105};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd125, 8'd130, 8'd107};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd106};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd106};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd125, 8'd132, 8'd106};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd106};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd106};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd123, 8'd127, 8'd104};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd126, 8'd126, 8'd105};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd123, 8'd126, 8'd105};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd122, 8'd123, 8'd105};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd123, 8'd125, 8'd105};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd121, 8'd127, 8'd104};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd105};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd104};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd125, 8'd128, 8'd105};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd108};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd129, 8'd125, 8'd108};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd129, 8'd124, 8'd107};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd131, 8'd125, 8'd109};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd134, 8'd127, 8'd111};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd131, 8'd128, 8'd113};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd132, 8'd129, 8'd116};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd128, 8'd129, 8'd115};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd112};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd127, 8'd130, 8'd115};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd128, 8'd130, 8'd115};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd127, 8'd135, 8'd112};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd127, 8'd134, 8'd114};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd127, 8'd134, 8'd113};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd127, 8'd134, 8'd113};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd114};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd114};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd123, 8'd131, 8'd112};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd111};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd124, 8'd131, 8'd113};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd112};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd111};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd114};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd114};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd130, 8'd133, 8'd114};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd129, 8'd134, 8'd113};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd130, 8'd135, 8'd115};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd132, 8'd138, 8'd115};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd133, 8'd142, 8'd117};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd133, 8'd143, 8'd117};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd130, 8'd140, 8'd115};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd128, 8'd138, 8'd114};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd113};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd112};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd111};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd112};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd127, 8'd135, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd129, 8'd138, 8'd114};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd134, 8'd143, 8'd115};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd138, 8'd146, 8'd122};
					endcase
				end
				`ybit'd29: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd113, 8'd121, 8'd110};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd116, 8'd124, 8'd113};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd115, 8'd125, 8'd108};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd114, 8'd129, 8'd107};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd115, 8'd128, 8'd107};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd116, 8'd126, 8'd109};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd113, 8'd124, 8'd107};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd111, 8'd122, 8'd105};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd109, 8'd124, 8'd103};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd107, 8'd125, 8'd103};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd109, 8'd127, 8'd105};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd111, 8'd129, 8'd105};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd113, 8'd128, 8'd105};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd113, 8'd128, 8'd108};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd113, 8'd128, 8'd109};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd116, 8'd126, 8'd110};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd120, 8'd126, 8'd116};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd122, 8'd128, 8'd115};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd110};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd117, 8'd131, 8'd106};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd112, 8'd127, 8'd104};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd102};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd111, 8'd123, 8'd103};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd115, 8'd123, 8'd109};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd118, 8'd126, 8'd115};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd123, 8'd126, 8'd116};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd124, 8'd127, 8'd116};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd124, 8'd128, 8'd111};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd111};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd119, 8'd128, 8'd108};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd117, 8'd126, 8'd106};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd114, 8'd124, 8'd103};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd112, 8'd124, 8'd101};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd98};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd109, 8'd122, 8'd95};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd108, 8'd118, 8'd92};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd108, 8'd118, 8'd94};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd109, 8'd119, 8'd95};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd98};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd112, 8'd124, 8'd102};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd104};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd115, 8'd125, 8'd101};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd99};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd111, 8'd121, 8'd96};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd113, 8'd123, 8'd99};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd115, 8'd125, 8'd100};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd118, 8'd128, 8'd109};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd115};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd133, 8'd139, 8'd131};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd133, 8'd139, 8'd131};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd134, 8'd135, 8'd130};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd133, 8'd129, 8'd126};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd131, 8'd126, 8'd123};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd129, 8'd123, 8'd120};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd128, 8'd123, 8'd119};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd125, 8'd121, 8'd117};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd125, 8'd120, 8'd117};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd127, 8'd122, 8'd120};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd130, 8'd125, 8'd127};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd131};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd129, 8'd129, 8'd129};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd125, 8'd125, 8'd125};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd125, 8'd127, 8'd115};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd128, 8'd129, 8'd114};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd112};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd115};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd131, 8'd128, 8'd119};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd131, 8'd128, 8'd121};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd134, 8'd128, 8'd123};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd123};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd137, 8'd129, 8'd119};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd138, 8'd126, 8'd115};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd136, 8'd124, 8'd111};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd133, 8'd121, 8'd109};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd106};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd133, 8'd121, 8'd109};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd130, 8'd120, 8'd108};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd129, 8'd120, 8'd108};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd127, 8'd119, 8'd106};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd126, 8'd118, 8'd105};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd124, 8'd120, 8'd103};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd104};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd127, 8'd124, 8'd107};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd134, 8'd123, 8'd109};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd131, 8'd122, 8'd107};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd129, 8'd118, 8'd106};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd129, 8'd119, 8'd106};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd127, 8'd120, 8'd104};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd105};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd123, 8'd127, 8'd104};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd106};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd104};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd105};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd124, 8'd135, 8'd105};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd124, 8'd136, 8'd106};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd121, 8'd134, 8'd104};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd103};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd121, 8'd133, 8'd103};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd105};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd125, 8'd129, 8'd104};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd125, 8'd129, 8'd106};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd123, 8'd129, 8'd105};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd105};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd105};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd121, 8'd126, 8'd103};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd122, 8'd126, 8'd103};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd122, 8'd127, 8'd103};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd121, 8'd129, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd121, 8'd129, 8'd103};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd121, 8'd129, 8'd103};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd120, 8'd129, 8'd101};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd103};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd103};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd124, 8'd127, 8'd105};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd106};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd108};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd106};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd129, 8'd122, 8'd106};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd132, 8'd125, 8'd109};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd130, 8'd126, 8'd111};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd129, 8'd126, 8'd111};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd124, 8'd125, 8'd111};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd122, 8'd124, 8'd110};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd123, 8'd125, 8'd111};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd123, 8'd124, 8'd110};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd110};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd124, 8'd127, 8'd111};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd110};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd110};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd125, 8'd130, 8'd110};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd124, 8'd128, 8'd111};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd121, 8'd125, 8'd108};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd121, 8'd125, 8'd108};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd121, 8'd128, 8'd110};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd110};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd110};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd111};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd111};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd112};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd126, 8'd131, 8'd111};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd126, 8'd131, 8'd111};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd129, 8'd134, 8'd111};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd113};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd129, 8'd138, 8'd113};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd136, 8'd111};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd125, 8'd135, 8'd111};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd111};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd111};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd110};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd111};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd109};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd110};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd128, 8'd137, 8'd108};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd130, 8'd138, 8'd114};
					endcase
				end
				`ybit'd30: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd107, 8'd118, 8'd101};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd107, 8'd122, 8'd103};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd108, 8'd123, 8'd103};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd109, 8'd124, 8'd101};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd111, 8'd127, 8'd101};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd111, 8'd127, 8'd101};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd110, 8'd125, 8'd106};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd110, 8'd121, 8'd104};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd108, 8'd120, 8'd100};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd105, 8'd122, 8'd99};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd107, 8'd125, 8'd100};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd109, 8'd125, 8'd99};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd108, 8'd124, 8'd101};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd106};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd106};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd116, 8'd122, 8'd112};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd117, 8'd123, 8'd112};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd118, 8'd126, 8'd112};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd119, 8'd128, 8'd106};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd114, 8'd127, 8'd101};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd97};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd110, 8'd120, 8'd96};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd111, 8'd119, 8'd102};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd111, 8'd117, 8'd106};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd115, 8'd121, 8'd110};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd117, 8'd123, 8'd112};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd120, 8'd126, 8'd113};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd120, 8'd127, 8'd106};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd116, 8'd128, 8'd104};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd104};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd113, 8'd125, 8'd103};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd111, 8'd122, 8'd101};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd110, 8'd121, 8'd99};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd94};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd108, 8'd121, 8'd93};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd106, 8'd119, 8'd91};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd108, 8'd118, 8'd93};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd108, 8'd118, 8'd93};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd109, 8'd120, 8'd95};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd98};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd113, 8'd126, 8'd99};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd113, 8'd126, 8'd100};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd97};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd97};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd110, 8'd120, 8'd96};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd111, 8'd122, 8'd98};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd116, 8'd128, 8'd104};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd120, 8'd132, 8'd112};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd125, 8'd136, 8'd118};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd129, 8'd136, 8'd128};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd129, 8'd135, 8'd132};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd130, 8'd132, 8'd129};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd127};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd125, 8'd124, 8'd128};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd125};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd125};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd125};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd125};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd132};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd125, 8'd125, 8'd135};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd129, 8'd129, 8'd140};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd127, 8'd129, 8'd136};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd122};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd125, 8'd127, 8'd116};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd124, 8'd125, 8'd109};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd108};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd108};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd114};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd130, 8'd124, 8'd121};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd130, 8'd125, 8'd119};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd132, 8'd127, 8'd120};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd137, 8'd126, 8'd116};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd136, 8'd124, 8'd112};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd106};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd106};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd107};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd133, 8'd120, 8'd108};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd130, 8'd121, 8'd109};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd128, 8'd121, 8'd108};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd126, 8'd120, 8'd106};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd104};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd125, 8'd119, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd127, 8'd120, 8'd107};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd134, 8'd120, 8'd109};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd107};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd107};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd107};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd130, 8'd122, 8'd106};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd128, 8'd124, 8'd105};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd124, 8'd125, 8'd103};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd126, 8'd127, 8'd104};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd103};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd106};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd121, 8'd133, 8'd105};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd123, 8'd136, 8'd101};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd101};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd105};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd106};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd105};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd126, 8'd129, 8'd105};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd124, 8'd127, 8'd102};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd122, 8'd128, 8'd102};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd103};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd105};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd106};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd122, 8'd128, 8'd104};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd120, 8'd129, 8'd104};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd121, 8'd132, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd120, 8'd131, 8'd102};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd122, 8'd132, 8'd105};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd102};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd120, 8'd129, 8'd100};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd121, 8'd129, 8'd101};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd106};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd127, 8'd128, 8'd106};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd128, 8'd126, 8'd105};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd104};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd107};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd129, 8'd125, 8'd106};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd108};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd110};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd109};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd108};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd107};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd107};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd108};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd121, 8'd122, 8'd108};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd108};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd108};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd109};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd122, 8'd123, 8'd109};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd120, 8'd121, 8'd108};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd120, 8'd122, 8'd108};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd122, 8'd127, 8'd106};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd123, 8'd130, 8'd107};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd123, 8'd131, 8'd108};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd110};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd111};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd126, 8'd131, 8'd109};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd109};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd109};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd108};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd126, 8'd134, 8'd110};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd125, 8'd133, 8'd109};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd108};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd124, 8'd131, 8'd109};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd111};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd111};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd110};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd123, 8'd133, 8'd109};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd123, 8'd133, 8'd110};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd109};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd109};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd109};
					endcase
				end
				`ybit'd31: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd105, 8'd117, 8'd95};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd103, 8'd118, 8'd93};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd103, 8'd119, 8'd94};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd104, 8'd119, 8'd96};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd106, 8'd122, 8'd96};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd108, 8'd124, 8'd98};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd108, 8'd123, 8'd103};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd107, 8'd118, 8'd101};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd105, 8'd117, 8'd97};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd102, 8'd119, 8'd95};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd103, 8'd121, 8'd97};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd104, 8'd120, 8'd94};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd109, 8'd120, 8'd99};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd113, 8'd119, 8'd107};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd113, 8'd120, 8'd108};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd114, 8'd120, 8'd110};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd115, 8'd121, 8'd109};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd117, 8'd126, 8'd107};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd115, 8'd125, 8'd100};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd97};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd107, 8'd120, 8'd94};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd107, 8'd117, 8'd93};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd107, 8'd116, 8'd98};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd107, 8'd114, 8'd97};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd109, 8'd116, 8'd100};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd114, 8'd121, 8'd104};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd117, 8'd124, 8'd107};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd117, 8'd129, 8'd106};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd117, 8'd129, 8'd105};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd113, 8'd125, 8'd103};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd100};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd109, 8'd121, 8'd99};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd108, 8'd120, 8'd98};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd95};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd109, 8'd122, 8'd94};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd106, 8'd120, 8'd92};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd106, 8'd116, 8'd91};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd106, 8'd116, 8'd91};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd108, 8'd119, 8'd93};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd98};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd114, 8'd127, 8'd101};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd115, 8'd128, 8'd102};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd114, 8'd127, 8'd101};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd97};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd110, 8'd120, 8'd96};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd109, 8'd121, 8'd97};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd102};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd120, 8'd132, 8'd112};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd122, 8'd132, 8'd120};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd132};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd138};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd121, 8'd126, 8'd137};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd121, 8'd123, 8'd137};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd118, 8'd120, 8'd136};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd117, 8'd120, 8'd136};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd116, 8'd118, 8'd138};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd116, 8'd117, 8'd140};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd116, 8'd117, 8'd140};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd146};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd119, 8'd121, 8'd151};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd122, 8'd125, 8'd149};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd125, 8'd127, 8'd141};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd123, 8'd127, 8'd126};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd122, 8'd124, 8'd113};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd122, 8'd123, 8'd107};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd106};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd106};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd111};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd126, 8'd121, 8'd117};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd127, 8'd122, 8'd117};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd130, 8'd125, 8'd118};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd135, 8'd124, 8'd114};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd133, 8'd121, 8'd109};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd106};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd127, 8'd115, 8'd103};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd127, 8'd115, 8'd103};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd128, 8'd116, 8'd104};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd127, 8'd115, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd127, 8'd115, 8'd103};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd129, 8'd117, 8'd105};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd133, 8'd119, 8'd108};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd131, 8'd117, 8'd106};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd128, 8'd116, 8'd104};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd124, 8'd115, 8'd102};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd125, 8'd114, 8'd102};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd106};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd107};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd133, 8'd119, 8'd108};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd107};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd108};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd133, 8'd119, 8'd106};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd131, 8'd122, 8'd105};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd128, 8'd124, 8'd106};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd125, 8'd122, 8'd104};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd124, 8'd120, 8'd103};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd122, 8'd123, 8'd102};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd122, 8'd129, 8'd103};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd101};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd127, 8'd137, 8'd103};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd127, 8'd136, 8'd107};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd105};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd120, 8'd130, 8'd103};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd120, 8'd129, 8'd102};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd119, 8'd130, 8'd103};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd121, 8'd132, 8'd104};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd99};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd103};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd102};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd102};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd102};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd121, 8'd132, 8'd102};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd100};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd103};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd101};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd101};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd101};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd101};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd124, 8'd128, 8'd104};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd124, 8'd128, 8'd105};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd124, 8'd128, 8'd105};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd127, 8'd127, 8'd107};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd105};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd108};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd108};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd105};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd105};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd105};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd106};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd119, 8'd120, 8'd106};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd106};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd107};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd107};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd119, 8'd120, 8'd106};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd116, 8'd118, 8'd104};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd118, 8'd120, 8'd106};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd120, 8'd125, 8'd105};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd120, 8'd128, 8'd105};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd107};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd123, 8'd131, 8'd108};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd105};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd105};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd104};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd104};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd106};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd123, 8'd131, 8'd107};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd106};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd105};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd104};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd122, 8'd132, 8'd107};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd120, 8'd130, 8'd106};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd121, 8'd131, 8'd106};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd124, 8'd134, 8'd106};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd122, 8'd133, 8'd105};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd124, 8'd131, 8'd108};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd107};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd120, 8'd128, 8'd105};
					endcase
				end
				`ybit'd32: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd103, 8'd115, 8'd92};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd101, 8'd117, 8'd90};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd101, 8'd117, 8'd90};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd101, 8'd118, 8'd91};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd103, 8'd119, 8'd93};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd104, 8'd120, 8'd94};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd104, 8'd120, 8'd94};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd103, 8'd118, 8'd95};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd103, 8'd115, 8'd93};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd103, 8'd115, 8'd91};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd104, 8'd115, 8'd91};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd105, 8'd117, 8'd93};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd108, 8'd116, 8'd96};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd112, 8'd117, 8'd103};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd114, 8'd118, 8'd105};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd115, 8'd118, 8'd109};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd113, 8'd120, 8'd105};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd111, 8'd123, 8'd102};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd96};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd108, 8'd121, 8'd93};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd104, 8'd117, 8'd91};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd105, 8'd114, 8'd93};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd103, 8'd112, 8'd91};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd104, 8'd112, 8'd91};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd105, 8'd115, 8'd97};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd109, 8'd118, 8'd101};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd114, 8'd123, 8'd105};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd116, 8'd130, 8'd107};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd105};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd115, 8'd127, 8'd103};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd111, 8'd123, 8'd99};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd102};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd99};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd112, 8'd125, 8'd96};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd110, 8'd123, 8'd95};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd111, 8'd120, 8'd93};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd107, 8'd115, 8'd92};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd108, 8'd116, 8'd93};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd110, 8'd118, 8'd95};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd111, 8'd126, 8'd100};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd114, 8'd131, 8'd100};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd116, 8'd133, 8'd102};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd114, 8'd130, 8'd104};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd112, 8'd124, 8'd101};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd110, 8'd119, 8'd99};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd109, 8'd120, 8'd103};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd113, 8'd125, 8'd107};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd116, 8'd130, 8'd115};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd116, 8'd129, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd116, 8'd126, 8'd138};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd116, 8'd124, 8'd147};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd115, 8'd122, 8'd152};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd114, 8'd118, 8'd150};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd113, 8'd117, 8'd149};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd112, 8'd116, 8'd149};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd112, 8'd115, 8'd154};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd112, 8'd115, 8'd156};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd111, 8'd113, 8'd153};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd111, 8'd112, 8'd159};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd113, 8'd116, 8'd158};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd115, 8'd121, 8'd156};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd119, 8'd123, 8'd142};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd117, 8'd124, 8'd123};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd119, 8'd122, 8'd110};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd119, 8'd121, 8'd109};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd120, 8'd121, 8'd106};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd111};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd116};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd118};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd125, 8'd119, 8'd115};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd128, 8'd123, 8'd113};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd130, 8'd123, 8'd108};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd106};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd125, 8'd114, 8'd102};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd124, 8'd114, 8'd102};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd124, 8'd114, 8'd102};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd126, 8'd114, 8'd102};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd126, 8'd113, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd126, 8'd113, 8'd104};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd128, 8'd115, 8'd106};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd107};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd107};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd130, 8'd116, 8'd105};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd127, 8'd115, 8'd103};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd126, 8'd113, 8'd104};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd125, 8'd112, 8'd103};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd127, 8'd114, 8'd105};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd130, 8'd116, 8'd105};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd130, 8'd116, 8'd105};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd130, 8'd116, 8'd105};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd106};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd105};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd133, 8'd119, 8'd106};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd105};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd128, 8'd117, 8'd102};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd122, 8'd115, 8'd99};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd100};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd123, 8'd124, 8'd101};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd100};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd126, 8'd136, 8'd102};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd130, 8'd137, 8'd103};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd127, 8'd137, 8'd102};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd124, 8'd134, 8'd100};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd120, 8'd129, 8'd100};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd119, 8'd128, 8'd101};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd121, 8'd129, 8'd100};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd124, 8'd132, 8'd103};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd126, 8'd136, 8'd102};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd102};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd102};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd102};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd125, 8'd135, 8'd101};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd103};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd103};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd126, 8'd135, 8'd106};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd128, 8'd134, 8'd106};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd129, 8'd133, 8'd107};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd107};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd105};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd105};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd125, 8'd129, 8'd107};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd122, 8'd125, 8'd104};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd120, 8'd121, 8'd107};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd105};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd103};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd103};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd118, 8'd119, 8'd104};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd118, 8'd120, 8'd101};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd119, 8'd121, 8'd105};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd119, 8'd121, 8'd105};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd104};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd105};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd116, 8'd118, 8'd102};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd117, 8'd119, 8'd103};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd118, 8'd123, 8'd103};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd118, 8'd127, 8'd103};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd123, 8'd128, 8'd105};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd123, 8'd131, 8'd107};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd106};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd106};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd105};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd103};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd103};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd121, 8'd130, 8'd103};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd103};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd121, 8'd131, 8'd104};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd104};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd122, 8'd132, 8'd104};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd132, 8'd104};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd124, 8'd135, 8'd105};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd125, 8'd135, 8'd106};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd123, 8'd133, 8'd106};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd121, 8'd131, 8'd104};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd120, 8'd125, 8'd104};
					endcase
				end
				`ybit'd33: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd100, 8'd113, 8'd86};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd98, 8'd113, 8'd87};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd87};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd99, 8'd116, 8'd84};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd101, 8'd118, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd102, 8'd118, 8'd92};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd102, 8'd118, 8'd92};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd101, 8'd116, 8'd93};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd101, 8'd113, 8'd92};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd101, 8'd114, 8'd90};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd101, 8'd113, 8'd89};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd100, 8'd112, 8'd88};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd105, 8'd114, 8'd94};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd110, 8'd114, 8'd100};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd112, 8'd116, 8'd102};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd112, 8'd115, 8'd106};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd110, 8'd118, 8'd103};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd108, 8'd120, 8'd98};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd108, 8'd121, 8'd94};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd105, 8'd118, 8'd90};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd103, 8'd116, 8'd90};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd102, 8'd111, 8'd90};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd101, 8'd110, 8'd89};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd102, 8'd110, 8'd89};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd102, 8'd112, 8'd88};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd106, 8'd116, 8'd92};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd113, 8'd123, 8'd99};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd115, 8'd131, 8'd104};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd117, 8'd133, 8'd106};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd116, 8'd129, 8'd104};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd103};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd113, 8'd125, 8'd105};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd103};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd115, 8'd128, 8'd100};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd114, 8'd126, 8'd99};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd95};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd108, 8'd116, 8'd93};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd109, 8'd117, 8'd94};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd111, 8'd120, 8'd96};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd112, 8'd126, 8'd100};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd115, 8'd131, 8'd105};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd106};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd115, 8'd129, 8'd111};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd112, 8'd123, 8'd110};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd109, 8'd117, 8'd107};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd108, 8'd117, 8'd113};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd110, 8'd120, 8'd115};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd112, 8'd123, 8'd127};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd134};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd112, 8'd118, 8'd150};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd112, 8'd116, 8'd159};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd110, 8'd114, 8'd163};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd108, 8'd114, 8'd167};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd107, 8'd113, 8'd165};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd107, 8'd113, 8'd165};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd106, 8'd112, 8'd163};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd106, 8'd112, 8'd165};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd106, 8'd111, 8'd166};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd105, 8'd109, 8'd170};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd106, 8'd111, 8'd166};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd109, 8'd113, 8'd159};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd111, 8'd116, 8'd151};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd111, 8'd120, 8'd134};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd113, 8'd120, 8'd120};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd112, 8'd118, 8'd114};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd114, 8'd117, 8'd116};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd114, 8'd116, 8'd122};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd114, 8'd114, 8'd127};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd124};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd117};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd113};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd127, 8'd119, 8'd104};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd123, 8'd116, 8'd102};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd123, 8'd114, 8'd101};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd122, 8'd112, 8'd100};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd121, 8'd111, 8'd99};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd123, 8'd111, 8'd99};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd120, 8'd113, 8'd102};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd120, 8'd113, 8'd102};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd126, 8'd113, 8'd104};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd132, 8'd118, 8'd106};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd131, 8'd117, 8'd106};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd129, 8'd115, 8'd104};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd125, 8'd114, 8'd101};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd124, 8'd111, 8'd102};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd124, 8'd111, 8'd102};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd125, 8'd113, 8'd103};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd129, 8'd114, 8'd103};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd129, 8'd115, 8'd104};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd129, 8'd115, 8'd104};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd128, 8'd114, 8'd104};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd128, 8'd114, 8'd101};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd128, 8'd114, 8'd101};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd126, 8'd114, 8'd100};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd124, 8'd112, 8'd99};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd121, 8'd108, 8'd99};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd118, 8'd110, 8'd100};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd123, 8'd118, 8'd100};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd100};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd133, 8'd101};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd102};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd126, 8'd136, 8'd102};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd122, 8'd132, 8'd99};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd119, 8'd128, 8'd100};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd117, 8'd126, 8'd99};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd119, 8'd128, 8'd99};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd101};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd125, 8'd135, 8'd101};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd128, 8'd135, 8'd102};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd129, 8'd136, 8'd103};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd136, 8'd103};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd127, 8'd134, 8'd102};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd126, 8'd136, 8'd102};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd123, 8'd133, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd104};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd125, 8'd134, 8'd105};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd127, 8'd136, 8'd107};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd132, 8'd141, 8'd112};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd136, 8'd142, 8'd114};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd138, 8'd142, 8'd117};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd136, 8'd140, 8'd115};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd135, 8'd139, 8'd114};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd132, 8'd136, 8'd111};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd106};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd125, 8'd129, 8'd103};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd123, 8'd124, 8'd104};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd100};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd116, 8'd119, 8'd98};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd114, 8'd118, 8'd97};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd115, 8'd117, 8'd97};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd114, 8'd121, 8'd97};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd116, 8'd122, 8'd99};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd116, 8'd122, 8'd99};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd118, 8'd121, 8'd100};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd118, 8'd121, 8'd100};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd116, 8'd119, 8'd97};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd116, 8'd119, 8'd98};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd115, 8'd120, 8'd101};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd120, 8'd122, 8'd102};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd122, 8'd127, 8'd104};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd105};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd122, 8'd130, 8'd106};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd107};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd107};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd126, 8'd130, 8'd105};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd104};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd122, 8'd131, 8'd104};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd123, 8'd132, 8'd105};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd124, 8'd133, 8'd106};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd125, 8'd135, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd125, 8'd136, 8'd102};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd127, 8'd138, 8'd103};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd137, 8'd103};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd128, 8'd139, 8'd105};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd127, 8'd138, 8'd104};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd126, 8'd137, 8'd106};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd123, 8'd134, 8'd103};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd120, 8'd125, 8'd104};
					endcase
				end
				`ybit'd34: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd97, 8'd113, 8'd84};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd96, 8'd112, 8'd83};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd85};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd85};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd100, 8'd117, 8'd84};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd100, 8'd117, 8'd84};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd100, 8'd116, 8'd90};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd99, 8'd115, 8'd88};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd87};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd96, 8'd112, 8'd85};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd96, 8'd112, 8'd85};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd99, 8'd111, 8'd87};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd103, 8'd112, 8'd92};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd105, 8'd113, 8'd95};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd105, 8'd113, 8'd95};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd106, 8'd114, 8'd96};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd106, 8'd118, 8'd98};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd107, 8'd119, 8'd96};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd107, 8'd120, 8'd90};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd105, 8'd118, 8'd90};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd102, 8'd115, 8'd89};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd102, 8'd112, 8'd90};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd99, 8'd108, 8'd88};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd100, 8'd109, 8'd90};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd102, 8'd111, 8'd90};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd104, 8'd116, 8'd94};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd112, 8'd124, 8'd102};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd113, 8'd132, 8'd104};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd114, 8'd133, 8'd105};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd114, 8'd132, 8'd106};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd113, 8'd131, 8'd105};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd106};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd106};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd104};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd116, 8'd131, 8'd102};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd114, 8'd124, 8'd98};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd111, 8'd117, 8'd99};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd109, 8'd115, 8'd101};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd111, 8'd117, 8'd103};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd110, 8'd122, 8'd110};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd111, 8'd127, 8'd114};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd112, 8'd127, 8'd119};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd110, 8'd124, 8'd123};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd108, 8'd119, 8'd123};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd106, 8'd112, 8'd124};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd103, 8'd111, 8'd126};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd106, 8'd114, 8'd134};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd107, 8'd114, 8'd140};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd105, 8'd113, 8'd148};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd106, 8'd111, 8'd158};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd108, 8'd110, 8'd165};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd108, 8'd110, 8'd167};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd107, 8'd109, 8'd168};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd105, 8'd110, 8'd168};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd105, 8'd110, 8'd168};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd104, 8'd109, 8'd167};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd104, 8'd109, 8'd167};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd104, 8'd108, 8'd168};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd103, 8'd107, 8'd168};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd103, 8'd108, 8'd167};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd103, 8'd108, 8'd162};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd103, 8'd110, 8'd155};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd104, 8'd112, 8'd141};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd108, 8'd113, 8'd131};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd107, 8'd112, 8'd127};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd108, 8'd113, 8'd128};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd108, 8'd111, 8'd135};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd107, 8'd110, 8'd136};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd107, 8'd110, 8'd134};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd112, 8'd113, 8'd123};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd100};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd120, 8'd115, 8'd101};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd123, 8'd113, 8'd101};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd121, 8'd111, 8'd99};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd98};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd100};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd121, 8'd112, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd120, 8'd111, 8'd102};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd125, 8'd114, 8'd105};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd129, 8'd116, 8'd107};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd130, 8'd116, 8'd105};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd127, 8'd113, 8'd102};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd125, 8'd111, 8'd100};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd124, 8'd111, 8'd102};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd122, 8'd109, 8'd100};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd123, 8'd111, 8'd101};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd127, 8'd112, 8'd103};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd127, 8'd113, 8'd104};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd127, 8'd113, 8'd102};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd126, 8'd112, 8'd101};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd124, 8'd110, 8'd99};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd122, 8'd109, 8'd100};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd121, 8'd108, 8'd99};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd118, 8'd106, 8'd97};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd113, 8'd103, 8'd94};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd117, 8'd106, 8'd97};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd120, 8'd114, 8'd100};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd99};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd127, 8'd104};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd102};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd127, 8'd130, 8'd103};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd124, 8'd127, 8'd101};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd122, 8'd125, 8'd98};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd120, 8'd124, 8'd101};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd121, 8'd126, 8'd99};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd124, 8'd129, 8'd101};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd127, 8'd130, 8'd100};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd128, 8'd131, 8'd102};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd129, 8'd132, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd132, 8'd103};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd129, 8'd132, 8'd102};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd128, 8'd133, 8'd103};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd100};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd100};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd99};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd125, 8'd130, 8'd102};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd129, 8'd133, 8'd106};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd135, 8'd139, 8'd112};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd145, 8'd148, 8'd121};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd151, 8'd153, 8'd127};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd152, 8'd155, 8'd128};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd151, 8'd154, 8'd127};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd149, 8'd152, 8'd125};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd142, 8'd147, 8'd120};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd137, 8'd141, 8'd114};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd131, 8'd135, 8'd109};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd125, 8'd129, 8'd104};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd121, 8'd123, 8'd101};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd118, 8'd120, 8'd100};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd116, 8'd117, 8'd98};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd115, 8'd118, 8'd97};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd115, 8'd119, 8'd97};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd115, 8'd119, 8'd97};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd115, 8'd120, 8'd97};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd116, 8'd121, 8'd99};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd115, 8'd120, 8'd98};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd115, 8'd118, 8'd97};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd114, 8'd116, 8'd95};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd117, 8'd119, 8'd98};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd120, 8'd122, 8'd101};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd125, 8'd127, 8'd106};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd128, 8'd130, 8'd109};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd131, 8'd133, 8'd112};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd134, 8'd136, 8'd114};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd135, 8'd138, 8'd116};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd133, 8'd136, 8'd113};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd132, 8'd134, 8'd112};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd130, 8'd135, 8'd112};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd132, 8'd136, 8'd111};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd132, 8'd138, 8'd112};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd133, 8'd141, 8'd114};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd136, 8'd145, 8'd116};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd140, 8'd149, 8'd116};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd139, 8'd149, 8'd115};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd136, 8'd147, 8'd113};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd136, 8'd147, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd136, 8'd147, 8'd113};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd132, 8'd142, 8'd109};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd124, 8'd128, 8'd106};
					endcase
				end
				`ybit'd35: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd95, 8'd111, 8'd82};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd96, 8'd111, 8'd82};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd97, 8'd112, 8'd83};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd100, 8'd116, 8'd86};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd100, 8'd117, 8'd82};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd100, 8'd117, 8'd81};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd100, 8'd116, 8'd85};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd98, 8'd113, 8'd83};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd96, 8'd111, 8'd84};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd94, 8'd110, 8'd83};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd94, 8'd110, 8'd83};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd97, 8'd109, 8'd84};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd101, 8'd111, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd100, 8'd111, 8'd88};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd99, 8'd112, 8'd88};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd100, 8'd114, 8'd90};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd102, 8'd116, 8'd91};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd104, 8'd118, 8'd92};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd106, 8'd120, 8'd90};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd104, 8'd119, 8'd90};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd103, 8'd117, 8'd90};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd101, 8'd112, 8'd89};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd99, 8'd109, 8'd88};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd100, 8'd109, 8'd90};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd101, 8'd110, 8'd91};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd104, 8'd117, 8'd96};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd102};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd112, 8'd131, 8'd103};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd115, 8'd133, 8'd106};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd115, 8'd132, 8'd107};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd114, 8'd132, 8'd106};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd115, 8'd132, 8'd107};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd116, 8'd133, 8'd107};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd107};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd114, 8'd129, 8'd105};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd113, 8'd123, 8'd103};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd111, 8'd116, 8'd105};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd108, 8'd111, 8'd109};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd109, 8'd112, 8'd113};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd107, 8'd116, 8'd122};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd106, 8'd119, 8'd127};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd107, 8'd119, 8'd135};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd106, 8'd116, 8'd140};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd105, 8'd113, 8'd141};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd102, 8'd108, 8'd142};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd102, 8'd107, 8'd146};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd103, 8'd108, 8'd151};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd103, 8'd108, 8'd156};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd102, 8'd108, 8'd161};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd164};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd168};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd105, 8'd106, 8'd169};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd105, 8'd106, 8'd170};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd103, 8'd107, 8'd170};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd103, 8'd107, 8'd170};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd102, 8'd106, 8'd169};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd102, 8'd106, 8'd166};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd168};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd100, 8'd105, 8'd161};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd100, 8'd106, 8'd155};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd101, 8'd107, 8'd147};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd100, 8'd106, 8'd143};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd101, 8'd108, 8'd145};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd101, 8'd107, 8'd148};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd101, 8'd107, 8'd148};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd103, 8'd108, 8'd142};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd108, 8'd112, 8'd126};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd112};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd102};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd121, 8'd115, 8'd101};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd122, 8'd112, 8'd100};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd99};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd119, 8'd109, 8'd97};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd119, 8'd109, 8'd98};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd120, 8'd112, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd121, 8'd114, 8'd107};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd124, 8'd115, 8'd106};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd128, 8'd115, 8'd106};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd129, 8'd115, 8'd105};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd125, 8'd111, 8'd101};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd124, 8'd110, 8'd100};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd122, 8'd109, 8'd100};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd120, 8'd108, 8'd99};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd121, 8'd109, 8'd100};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd122, 8'd111, 8'd101};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd124, 8'd110, 8'd101};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd126, 8'd112, 8'd101};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd125, 8'd111, 8'd99};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd121, 8'd108, 8'd97};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd117, 8'd104, 8'd96};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd116, 8'd104, 8'd94};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd112, 8'd101, 8'd92};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd110, 8'd101, 8'd93};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd112, 8'd102, 8'd93};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd118, 8'd109, 8'd99};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd124, 8'd115, 8'd99};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd127, 8'd121, 8'd103};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd130, 8'd126, 8'd103};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd129, 8'd125, 8'd104};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd102};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd126, 8'd122, 8'd103};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd124, 8'd123, 8'd101};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd124, 8'd123, 8'd102};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd127, 8'd124, 8'd104};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd128, 8'd124, 8'd103};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd129, 8'd125, 8'd102};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd126, 8'd102};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd102};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd103};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd128, 8'd126, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd101};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd102};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd127, 8'd127, 8'd100};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd130, 8'd130, 8'd104};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd114};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd129};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd164, 8'd162, 8'd138};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd167, 8'd165, 8'd141};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd166, 8'd164, 8'd140};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd164, 8'd162, 8'd138};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd158, 8'd157, 8'd131};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd145, 8'd148, 8'd120};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd134, 8'd138, 8'd110};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd125, 8'd131, 8'd100};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd122, 8'd126, 8'd99};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd119, 8'd121, 8'd98};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd116, 8'd119, 8'd96};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd114, 8'd116, 8'd95};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd115, 8'd116, 8'd95};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd113, 8'd116, 8'd94};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd112, 8'd116, 8'd95};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd113, 8'd117, 8'd96};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd113, 8'd117, 8'd96};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd113, 8'd116, 8'd95};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd114, 8'd117, 8'd96};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd117, 8'd119, 8'd99};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd106};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd132, 8'd129, 8'd111};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd116};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd118};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd122};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd124};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd125};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd122};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd120};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd144, 8'd143, 8'd121};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd146, 8'd146, 8'd123};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd145, 8'd149, 8'd125};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd151, 8'd154, 8'd128};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd155, 8'd160, 8'd128};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd155, 8'd160, 8'd128};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd153, 8'd160, 8'd127};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd154, 8'd160, 8'd128};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd152, 8'd158, 8'd127};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd146, 8'd153, 8'd122};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd137, 8'd141, 8'd118};
					endcase
				end
				`ybit'd36: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd93, 8'd109, 8'd80};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd96, 8'd110, 8'd82};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd99, 8'd112, 8'd84};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd99, 8'd116, 8'd84};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd99, 8'd116, 8'd84};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd97, 8'd114, 8'd82};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd97, 8'd114, 8'd82};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd99, 8'd112, 8'd84};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd96, 8'd109, 8'd83};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd92, 8'd107, 8'd80};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd91, 8'd107, 8'd80};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd94, 8'd107, 8'd81};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd95, 8'd109, 8'd84};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd97, 8'd111, 8'd83};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd97, 8'd112, 8'd84};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd97, 8'd113, 8'd85};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd99, 8'd115, 8'd89};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd103, 8'd119, 8'd93};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd105, 8'd120, 8'd95};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd104, 8'd119, 8'd97};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd103, 8'd118, 8'd98};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd103, 8'd114, 8'd97};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd99, 8'd110, 8'd94};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd101, 8'd109, 8'd98};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd100, 8'd110, 8'd101};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd102, 8'd115, 8'd106};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd108, 8'd121, 8'd111};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd109, 8'd125, 8'd114};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd111, 8'd127, 8'd116};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd111, 8'd126, 8'd117};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd111, 8'd126, 8'd118};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd110, 8'd125, 8'd119};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd110, 8'd125, 8'd119};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd112, 8'd125, 8'd119};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd118};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd108, 8'd120, 8'd118};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd109, 8'd113, 8'd123};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd106, 8'd109, 8'd126};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd104, 8'd108, 8'd132};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd102, 8'd109, 8'd138};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd101, 8'd109, 8'd143};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd102, 8'd110, 8'd148};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd102, 8'd109, 8'd153};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd102, 8'd108, 8'd156};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd156};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd101, 8'd104, 8'd157};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd159};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd101, 8'd105, 8'd163};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd165};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd166};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd101, 8'd104, 8'd167};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd167};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd167};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd97, 8'd102, 8'd158};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd97, 8'd102, 8'd156};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd97, 8'd104, 8'd149};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd99, 8'd105, 8'd151};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd99, 8'd106, 8'd145};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd100, 8'd107, 8'd146};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd102, 8'd110, 8'd140};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd109, 8'd113, 8'd123};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd116, 8'd117, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd121, 8'd115, 8'd102};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd122, 8'd112, 8'd100};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd121, 8'd111, 8'd100};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd118, 8'd108, 8'd97};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd117, 8'd107, 8'd95};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd117, 8'd110, 8'd98};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd118, 8'd115, 8'd110};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd122, 8'd117, 8'd108};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd126, 8'd115, 8'd105};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd127, 8'd114, 8'd105};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd126, 8'd113, 8'd104};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd122, 8'd109, 8'd100};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd119, 8'd106, 8'd97};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd117, 8'd108, 8'd99};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd118, 8'd108, 8'd99};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd103};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd122, 8'd113, 8'd105};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd122, 8'd113, 8'd103};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd100};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd117, 8'd104, 8'd95};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd114, 8'd101, 8'd93};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd111, 8'd101, 8'd92};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd109, 8'd99, 8'd90};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd107, 8'd98, 8'd93};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd110, 8'd100, 8'd91};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd119, 8'd106, 8'd97};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd123, 8'd111, 8'd95};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd116, 8'd102};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd103};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd131, 8'd119, 8'd103};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd131, 8'd118, 8'd103};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd102};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd128, 8'd119, 8'd102};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd129, 8'd120, 8'd102};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd129, 8'd120, 8'd103};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd129, 8'd120, 8'd103};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd131, 8'd120, 8'd101};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd129, 8'd121, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd122, 8'd102};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd130, 8'd123, 8'd103};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd130, 8'd122, 8'd103};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd129, 8'd122, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd129, 8'd122, 8'd102};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd129, 8'd121, 8'd102};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd129, 8'd122, 8'd102};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd131, 8'd125, 8'd105};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd167, 8'd165, 8'd142};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd171, 8'd169, 8'd146};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd171, 8'd169, 8'd146};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd169, 8'd167, 8'd144};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd162, 8'd162, 8'd137};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd124};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd110};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd125, 8'd126, 8'd101};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd121, 8'd122, 8'd98};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd98};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd96};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd95};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd115, 8'd112, 8'd93};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd111, 8'd113, 8'd94};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd110, 8'd112, 8'd94};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd109, 8'd112, 8'd93};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd109, 8'd112, 8'd93};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd109, 8'd112, 8'd91};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd112, 8'd115, 8'd94};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd120, 8'd121, 8'd103};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd110};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd139, 8'd136, 8'd118};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd122};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd148, 8'd145, 8'd126};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd152, 8'd149, 8'd130};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd132};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd131};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd128};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd146, 8'd126};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd148, 8'd147, 8'd126};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd152, 8'd151, 8'd130};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd158, 8'd157, 8'd136};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd163, 8'd162, 8'd138};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd167, 8'd168, 8'd141};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd167, 8'd168, 8'd141};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd165, 8'd166, 8'd137};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd165, 8'd166, 8'd139};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd164, 8'd165, 8'd138};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd159, 8'd161, 8'd134};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd153, 8'd154, 8'd129};
					endcase
				end
				`ybit'd37: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd92, 8'd111, 8'd81};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd95, 8'd112, 8'd77};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd96, 8'd112, 8'd78};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd95, 8'd113, 8'd81};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd96, 8'd113, 8'd81};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd97, 8'd111, 8'd83};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd97, 8'd111, 8'd84};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd99, 8'd109, 8'd84};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd95, 8'd108, 8'd82};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd91, 8'd104, 8'd78};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd91, 8'd104, 8'd78};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd92, 8'd105, 8'd79};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd93, 8'd109, 8'd80};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd93, 8'd110, 8'd80};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd94, 8'd110, 8'd81};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd96, 8'd112, 8'd83};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd97, 8'd116, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd100, 8'd118, 8'd91};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd102, 8'd118, 8'd103};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd102, 8'd118, 8'd107};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd102, 8'd118, 8'd108};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd101, 8'd114, 8'd105};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd98, 8'd110, 8'd106};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd98, 8'd109, 8'd110};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd99, 8'd109, 8'd114};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd101, 8'd113, 8'd120};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd104, 8'd117, 8'd124};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd105, 8'd118, 8'd129};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd105, 8'd117, 8'd129};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd106, 8'd118, 8'd133};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd106, 8'd118, 8'd134};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd105, 8'd116, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd105, 8'd116, 8'd136};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd105, 8'd116, 8'd135};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd104, 8'd115, 8'd134};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd104, 8'd112, 8'd137};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd102, 8'd111, 8'd139};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd99, 8'd107, 8'd142};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd99, 8'd105, 8'd146};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd101, 8'd104, 8'd153};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd100, 8'd105, 8'd158};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd99, 8'd105, 8'd160};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd161};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd162};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd166};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd100, 8'd103, 8'd166};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd101, 8'd105, 8'd168};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd167};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd100, 8'd103, 8'd166};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd95, 8'd100, 8'd163};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd163};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd162};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd162};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd162};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd163};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd158};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd153};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd98, 8'd104, 8'd152};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd98, 8'd106, 8'd143};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd100, 8'd110, 8'd132};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd101, 8'd110, 8'd127};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd104, 8'd112, 8'd124};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd111, 8'd114, 8'd116};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd108};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd121, 8'd113, 8'd100};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd121, 8'd111, 8'd99};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd118, 8'd110, 8'd97};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd115, 8'd107, 8'd94};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd116, 8'd108, 8'd93};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd116, 8'd110, 8'd95};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd111};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd121, 8'd115, 8'd111};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd127, 8'd117, 8'd107};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd128, 8'd115, 8'd106};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd124, 8'd111, 8'd102};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd121, 8'd108, 8'd99};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd117, 8'd107, 8'd98};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd118, 8'd107, 8'd97};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd117, 8'd111, 8'd106};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd121, 8'd114, 8'd108};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd120, 8'd113, 8'd107};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd119, 8'd112, 8'd105};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd116, 8'd108, 8'd102};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd113, 8'd103, 8'd96};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd109, 8'd98, 8'd94};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd108, 8'd99, 8'd94};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd106, 8'd97, 8'd91};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd103, 8'd98, 8'd92};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd108, 8'd100, 8'd92};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd119, 8'd105, 8'd94};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd124, 8'd109, 8'd98};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd130, 8'd114, 8'd101};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd131, 8'd115, 8'd103};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd134, 8'd117, 8'd103};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd103};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd102};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd133, 8'd118, 8'd104};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd134, 8'd118, 8'd105};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd134, 8'd119, 8'd105};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd132, 8'd117, 8'd103};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd132, 8'd116, 8'd103};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd133, 8'd116, 8'd103};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd133, 8'd116, 8'd103};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd132, 8'd117, 8'd102};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd104};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd130, 8'd118, 8'd102};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd132, 8'd117, 8'd103};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd132, 8'd117, 8'd104};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd136, 8'd122, 8'd106};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd145, 8'd137, 8'd120};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd159, 8'd152, 8'd133};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd168, 8'd162, 8'd142};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd170, 8'd163, 8'd144};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd170, 8'd164, 8'd144};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd170, 8'd164, 8'd140};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd163, 8'd157, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd148, 8'd142, 8'd121};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd131, 8'd126, 8'd105};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd98};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd97};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd118, 8'd115, 8'd96};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd95};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd117, 8'd112, 8'd95};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd117, 8'd110, 8'd94};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd115, 8'd110, 8'd93};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd108, 8'd110, 8'd92};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd88};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd105, 8'd106, 8'd90};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd106, 8'd108, 8'd91};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd111, 8'd113, 8'd96};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd120, 8'd121, 8'd103};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd142, 8'd139, 8'd122};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd126};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd151, 8'd148, 8'd129};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd133};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd135};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd133};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd149, 8'd146, 8'd128};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd124};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd126};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd130};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd158, 8'd155, 8'd136};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd165, 8'd162, 8'd141};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd168, 8'd166, 8'd142};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd168, 8'd166, 8'd141};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd165, 8'd163, 8'd137};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd164, 8'd162, 8'd137};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd163, 8'd163, 8'd136};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd162, 8'd162, 8'd136};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd162, 8'd160, 8'd133};
					endcase
				end
				`ybit'd38: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd92, 8'd112, 8'd75};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd95, 8'd112, 8'd76};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd94, 8'd112, 8'd76};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd92, 8'd111, 8'd79};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd93, 8'd110, 8'd78};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd94, 8'd107, 8'd81};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd94, 8'd107, 8'd81};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd96, 8'd106, 8'd81};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd94, 8'd107, 8'd81};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd92, 8'd105, 8'd79};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd90, 8'd103, 8'd77};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd91, 8'd104, 8'd78};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd92, 8'd108, 8'd79};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd91, 8'd107, 8'd78};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd94, 8'd110, 8'd81};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd94, 8'd110, 8'd81};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd96, 8'd114, 8'd88};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd97};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd100, 8'd115, 8'd111};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd101, 8'd115, 8'd118};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd101, 8'd114, 8'd123};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd101, 8'd111, 8'd119};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd99, 8'd108, 8'd122};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd98, 8'd106, 8'd126};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd99, 8'd107, 8'd131};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd100, 8'd108, 8'd139};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd102, 8'd110, 8'd142};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd101, 8'd109, 8'd145};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd102, 8'd109, 8'd149};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd102, 8'd109, 8'd149};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd102, 8'd109, 8'd150};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd101, 8'd108, 8'd152};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd102, 8'd108, 8'd152};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd100, 8'd107, 8'd151};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd102, 8'd108, 8'd152};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd102, 8'd107, 8'd152};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd100, 8'd106, 8'd153};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd156};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd101, 8'd103, 8'd162};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd98, 8'd103, 8'd161};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd164};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd164};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd162};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd167};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd162};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd93, 8'd99, 8'd161};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd93, 8'd99, 8'd161};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd93, 8'd99, 8'd161};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd93, 8'd99, 8'd161};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd94, 8'd99, 8'd158};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd95, 8'd101, 8'd152};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd96, 8'd103, 8'd143};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd101, 8'd105, 8'd136};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd103, 8'd109, 8'd128};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd104, 8'd112, 8'd117};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd107, 8'd113, 8'd112};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd107, 8'd113, 8'd109};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd110, 8'd114, 8'd104};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd98};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd118, 8'd110, 8'd97};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd118, 8'd108, 8'd96};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd116, 8'd108, 8'd95};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd114, 8'd106, 8'd93};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd116, 8'd109, 8'd93};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd95};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd112};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd121, 8'd117, 8'd112};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd124, 8'd118, 8'd113};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd124, 8'd116, 8'd109};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd122, 8'd113, 8'd106};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd118, 8'd109, 8'd103};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd114, 8'd109, 8'd104};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd116, 8'd110, 8'd103};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd113};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd120, 8'd116, 8'd113};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd117, 8'd113, 8'd111};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd107};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd111, 8'd107, 8'd104};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd107, 8'd103, 8'd100};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd107, 8'd101, 8'd95};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd108, 8'd100, 8'd94};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd107, 8'd99, 8'd93};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd103, 8'd98, 8'd92};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd109, 8'd101, 8'd93};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd118, 8'd104, 8'd93};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd124, 8'd109, 8'd98};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd131, 8'd115, 8'd102};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd132, 8'd116, 8'd101};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd132, 8'd116, 8'd101};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd102};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd104};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd104};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd104};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd133, 8'd117, 8'd104};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd131, 8'd115, 8'd102};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd101};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd132, 8'd114, 8'd101};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd132, 8'd116, 8'd101};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd134, 8'd116, 8'd104};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd134, 8'd116, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd133, 8'd115, 8'd101};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd132, 8'd116, 8'd103};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd131, 8'd115, 8'd102};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd136, 8'd121, 8'd106};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd144, 8'd136, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd157, 8'd150, 8'd131};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd164, 8'd157, 8'd138};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd164, 8'd157, 8'd138};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd163, 8'd156, 8'd138};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd161, 8'd154, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd154, 8'd147, 8'd130};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd139, 8'd132, 8'd115};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd125, 8'd118, 8'd102};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd98};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd98};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd98};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd98};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd122, 8'd111, 8'd97};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd118, 8'd111, 8'd95};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd116, 8'd110, 8'd94};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd107, 8'd109, 8'd91};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd106, 8'd109, 8'd90};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd105, 8'd106, 8'd90};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd90};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd95};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd103};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd141, 8'd139, 8'd122};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd126};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd151, 8'd148, 8'd129};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd133};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd133};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd151, 8'd148, 8'd129};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd123};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd120};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd120};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd126};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd153, 8'd150, 8'd131};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd137};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd162, 8'd159, 8'd140};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd137};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd132};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd153, 8'd150, 8'd130};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd133};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd155, 8'd154, 8'd133};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
					endcase
				end
				`ybit'd39: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd92, 8'd112, 8'd75};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd91, 8'd111, 8'd74};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd90, 8'd110, 8'd74};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd91, 8'd108, 8'd76};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd89, 8'd106, 8'd73};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd90, 8'd104, 8'd77};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd91, 8'd103, 8'd77};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd93, 8'd103, 8'd78};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd94, 8'd104, 8'd79};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd91, 8'd104, 8'd78};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd89, 8'd102, 8'd76};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd90, 8'd103, 8'd77};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd87, 8'd103, 8'd74};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd91, 8'd107, 8'd78};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd91, 8'd108, 8'd78};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd91, 8'd110, 8'd78};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd95, 8'd113, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd96, 8'd114, 8'd96};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd96, 8'd110, 8'd113};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd98, 8'd110, 8'd125};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd98, 8'd110, 8'd125};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd96, 8'd107, 8'd126};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd94, 8'd104, 8'd129};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd96, 8'd103, 8'd133};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd96, 8'd104, 8'd143};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd98, 8'd105, 8'd151};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd157};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd155};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd159};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd99, 8'd104, 8'd160};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd98, 8'd103, 8'd160};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd98, 8'd103, 8'd161};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd99, 8'd102, 8'd165};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd97, 8'd102, 8'd164};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd166};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd163};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd95, 8'd101, 8'd163};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd95, 8'd98, 8'd163};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd162};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd161};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd91, 8'd97, 8'd161};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd162};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd91, 8'd99, 8'd162};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd162};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd161};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd161};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd162};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd154};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd97, 8'd104, 8'd144};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd102, 8'd106, 8'd128};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd102, 8'd110, 8'd120};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd106, 8'd109, 8'd113};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd107, 8'd112, 8'd107};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd106, 8'd113, 8'd103};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd111, 8'd113, 8'd99};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd109, 8'd115, 8'd95};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd95};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd116, 8'd109, 8'd93};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd92};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd92};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd90};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd93};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd114, 8'd115, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd109};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd116};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd116};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd125, 8'd119, 8'd114};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd121, 8'd115, 8'd109};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd117, 8'd110, 8'd105};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd115, 8'd108, 8'd103};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd117, 8'd116, 8'd111};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd117};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd114};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd109};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd107};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd104};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd102};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd109, 8'd104, 8'd101};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd107, 8'd102, 8'd99};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd94};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd109, 8'd100, 8'd93};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd116, 8'd105, 8'd96};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd126, 8'd108, 8'd94};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd112, 8'd99};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd129, 8'd113, 8'd100};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd131, 8'd112, 8'd101};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd100};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd132, 8'd114, 8'd100};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd133, 8'd115, 8'd103};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd133, 8'd115, 8'd103};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd132, 8'd114, 8'd101};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd98};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd98};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd99};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd100};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd132, 8'd114, 8'd100};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd132, 8'd114, 8'd100};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd133, 8'd115, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd132, 8'd114, 8'd102};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd100};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd129, 8'd113, 8'd100};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd134, 8'd119, 8'd106};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd142, 8'd135, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd155, 8'd148, 8'd130};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd156, 8'd153, 8'd134};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd158, 8'd152, 8'd133};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd156, 8'd149, 8'd131};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd154, 8'd147, 8'd129};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd147, 8'd140, 8'd124};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd135, 8'd128, 8'd112};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd126, 8'd119, 8'd103};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd121, 8'd114, 8'd98};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd120, 8'd112, 8'd99};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd122, 8'd112, 8'd100};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd124, 8'd114, 8'd101};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd123, 8'd114, 8'd99};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd123, 8'd116, 8'd98};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd119, 8'd114, 8'd95};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd111, 8'd113, 8'd92};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd107, 8'd110, 8'd88};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd105, 8'd107, 8'd89};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd90};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd113, 8'd109, 8'd95};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd124, 8'd116, 8'd100};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd110};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd137, 8'd135, 8'd116};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd140, 8'd140, 8'd119};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd145, 8'd144, 8'd124};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd148, 8'd145, 8'd126};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd146, 8'd143, 8'd126};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd121};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd136, 8'd133, 8'd118};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd133, 8'd131, 8'd116};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd137, 8'd135, 8'd120};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd142, 8'd139, 8'd124};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd150, 8'd147, 8'd130};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd154, 8'd151, 8'd132};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd151, 8'd148, 8'd132};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd127};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd142, 8'd141, 8'd123};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd140, 8'd139, 8'd121};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd123};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd147, 8'd144, 8'd126};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd128};
					endcase
				end
				`ybit'd40: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd91, 8'd111, 8'd73};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd89, 8'd109, 8'd72};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd87, 8'd107, 8'd70};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd88, 8'd105, 8'd73};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd88, 8'd104, 8'd76};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd88, 8'd101, 8'd75};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd89, 8'd102, 8'd75};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd90, 8'd100, 8'd75};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd90, 8'd100, 8'd75};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd89, 8'd102, 8'd76};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd89, 8'd102, 8'd76};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd89, 8'd102, 8'd76};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd88, 8'd104, 8'd75};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd87, 8'd103, 8'd74};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd90, 8'd107, 8'd77};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd90, 8'd109, 8'd77};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd93, 8'd112, 8'd78};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd94, 8'd112, 8'd89};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd94, 8'd109, 8'd106};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd94, 8'd107, 8'd117};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd94, 8'd106, 8'd121};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd94, 8'd105, 8'd123};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd92, 8'd102, 8'd127};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd136};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd95, 8'd102, 8'd147};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd158};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd97, 8'd100, 8'd164};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd97, 8'd100, 8'd163};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd162};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd164};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd165};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd165};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd94, 8'd99, 8'd161};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd92, 8'd99, 8'd161};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd160};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd161};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd161};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd91, 8'd98, 8'd155};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd94, 8'd101, 8'd147};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd96, 8'd105, 8'd133};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd103, 8'd108, 8'd117};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd106, 8'd111, 8'd104};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd105, 8'd110, 8'd99};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd105, 8'd112, 8'd93};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd108, 8'd110, 8'd90};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd107, 8'd110, 8'd90};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd107, 8'd113, 8'd93};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd111, 8'd111, 8'd93};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd91};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd114, 8'd107, 8'd91};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd92};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd91};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd91};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd94};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd114, 8'd115, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd111};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd115};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd122};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd119};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd114};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd114, 8'd112, 8'd110};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd108};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd110};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd115};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd116, 8'd116, 8'd116};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd111};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd111};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd110};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd115, 8'd111, 8'd108};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd116, 8'd110, 8'd107};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd112, 8'd107, 8'd105};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd108, 8'd103, 8'd98};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd95};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd117, 8'd105, 8'd96};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd126, 8'd108, 8'd94};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd97};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd128, 8'd112, 8'd99};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd100};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd100};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd99};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd101};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd101};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd101};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd130, 8'd112, 8'd98};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd128, 8'd110, 8'd96};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd129, 8'd111, 8'd99};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd111, 8'd99};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd99};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd99};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd100};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd101};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd129, 8'd111, 8'd99};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd128, 8'd112, 8'd99};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd132, 8'd117, 8'd104};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd139, 8'd132, 8'd116};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd153, 8'd146, 8'd128};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd154, 8'd151, 8'd133};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd156, 8'd149, 8'd131};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd154, 8'd147, 8'd129};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd152, 8'd145, 8'd127};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd148, 8'd141, 8'd125};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd140, 8'd133, 8'd117};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd135, 8'd128, 8'd112};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd132, 8'd125, 8'd109};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd132, 8'd124, 8'd111};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd133, 8'd123, 8'd111};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd134, 8'd124, 8'd112};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd135, 8'd126, 8'd111};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd132, 8'd125, 8'd107};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd127, 8'd123, 8'd104};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd114, 8'd116, 8'd96};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd108, 8'd111, 8'd90};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd110, 8'd106, 8'd89};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd113, 8'd103, 8'd91};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd114, 8'd105, 8'd92};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd119, 8'd112, 8'd96};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd124, 8'd121, 8'd104};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd128, 8'd127, 8'd107};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd112};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd115};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd115};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd133, 8'd130, 8'd112};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd108};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd108};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd110};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd132, 8'd129, 8'd114};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd121};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd145, 8'd142, 8'd125};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd147, 8'd144, 8'd125};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd123};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd117};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd136, 8'd133, 8'd116};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd120};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd124};
					endcase
				end
				`ybit'd41: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd87, 8'd106, 8'd74};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd88, 8'd105, 8'd75};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd73};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd87, 8'd103, 8'd76};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd75};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd86, 8'd98, 8'd74};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd85, 8'd97, 8'd73};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd85, 8'd97, 8'd73};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd86, 8'd99, 8'd73};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd87, 8'd102, 8'd74};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd87, 8'd103, 8'd76};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd89, 8'd106, 8'd76};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd89, 8'd108, 8'd76};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd92, 8'd112, 8'd77};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd90, 8'd109, 8'd83};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd90, 8'd107, 8'd95};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd91, 8'd106, 8'd101};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd91, 8'd105, 8'd106};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd92, 8'd102, 8'd111};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd92, 8'd101, 8'd116};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd91, 8'd99, 8'd128};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd93, 8'd100, 8'd141};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd154};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd161};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd163};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd163};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd163};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd164};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd161};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd160};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd160};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd160};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd88, 8'd96, 8'd160};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd159};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd161};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd161};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd156};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd95, 8'd102, 8'd146};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd97, 8'd107, 8'd132};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd101, 8'd108, 8'd113};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd103, 8'd111, 8'd103};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd105, 8'd109, 8'd93};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd106, 8'd110, 8'd89};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd105, 8'd108, 8'd87};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd106, 8'd109, 8'd88};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd108, 8'd111, 8'd90};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd108, 8'd111, 8'd90};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd87};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd90};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd89};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd89};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd89};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd114, 8'd110, 8'd94};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd103};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd109};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd116};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd120};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd120};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd117};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd109, 8'd109, 8'd109};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd111, 8'd111, 8'd111};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd116};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd117};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd117};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd120, 8'd116, 8'd113};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd119, 8'd114, 8'd110};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd116, 8'd112, 8'd108};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd112, 8'd107, 8'd101};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd112, 8'd103, 8'd96};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd119, 8'd104, 8'd93};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd122, 8'd109, 8'd97};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd125, 8'd109, 8'd96};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd97};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd97};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd97};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd97};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd96};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd129, 8'd113, 8'd100};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd129, 8'd113, 8'd98};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd128, 8'd110, 8'd96};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd128, 8'd110, 8'd96};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd129, 8'd116, 8'd103};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd140, 8'd134, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd155, 8'd148, 8'd129};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd133};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd133};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd132};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd156, 8'd149, 8'd131};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd154, 8'd147, 8'd129};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd150, 8'd143, 8'd125};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd149, 8'd142, 8'd123};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd147, 8'd139, 8'd121};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd145, 8'd138, 8'd120};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd146, 8'd139, 8'd122};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd147, 8'd140, 8'd123};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd149, 8'd141, 8'd123};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd121};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd136, 8'd134, 8'd113};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd100};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd93};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd89};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd90};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd89};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd115, 8'd107, 8'd94};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd97};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd99};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd123, 8'd122, 8'd102};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd124, 8'd123, 8'd103};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd101};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd117, 8'd113, 8'd101};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd115, 8'd111, 8'd99};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd116, 8'd112, 8'd100};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd119, 8'd115, 8'd103};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd130, 8'd124, 8'd108};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd138, 8'd131, 8'd115};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd142, 8'd135, 8'd119};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd117};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd133, 8'd130, 8'd115};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd112};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd112};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd112};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd133, 8'd133, 8'd114};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd118};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd119};
					endcase
				end
				`ybit'd42: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd84, 8'd103, 8'd71};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd85, 8'd102, 8'd72};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd74};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd74};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd85, 8'd97, 8'd73};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd82, 8'd95, 8'd70};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd82, 8'd94, 8'd70};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd83, 8'd96, 8'd70};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd74};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd73};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd89, 8'd105, 8'd75};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd90, 8'd109, 8'd77};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd90, 8'd109, 8'd76};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd88, 8'd107, 8'd73};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd87, 8'd105, 8'd81};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd89, 8'd105, 8'd87};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd90, 8'd105, 8'd91};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd91, 8'd103, 8'd98};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd90, 8'd100, 8'd103};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd90, 8'd99, 8'd115};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd90, 8'd99, 8'd129};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd147};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd95, 8'd100, 8'd154};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd95, 8'd100, 8'd155};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd156};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd156};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd95, 8'd100, 8'd156};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd95, 8'd100, 8'd158};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd160};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd163};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd161};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd160};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd161};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd157};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd157};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd158};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd157};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd88, 8'd97, 8'd156};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd158};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd159};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd159};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd158};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd87, 8'd95, 8'd158};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd160};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd160};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd93, 8'd98, 8'd156};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd93, 8'd100, 8'd145};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd96, 8'd105, 8'd132};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd98, 8'd105, 8'd116};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd100, 8'd107, 8'd105};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd104, 8'd109, 8'd93};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd105, 8'd109, 8'd88};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd105, 8'd108, 8'd87};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd86};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd86};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd106, 8'd109, 8'd88};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd86};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd87};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd85};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd86};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd88};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd116, 8'd106, 8'd93};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd102};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd109};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd114};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd118, 8'd118, 8'd118};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd119};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd114, 8'd114, 8'd114};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd114, 8'd114, 8'd114};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd117, 8'd116, 8'd116};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd118};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd117};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd117, 8'd113, 8'd110};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd119, 8'd111, 8'd104};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd117, 8'd107, 8'd100};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd114, 8'd103, 8'd99};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd112, 8'd102, 8'd95};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd116, 8'd102, 8'd92};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd118, 8'd104, 8'd93};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd121, 8'd105, 8'd92};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd121, 8'd105, 8'd92};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd121, 8'd105, 8'd92};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd123, 8'd107, 8'd94};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd123, 8'd107, 8'd94};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd123, 8'd106, 8'd97};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd123, 8'd106, 8'd97};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd123, 8'd106, 8'd97};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd123, 8'd108, 8'd95};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd125, 8'd109, 8'd96};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd96};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd127, 8'd108, 8'd95};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd126, 8'd109, 8'd95};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd125, 8'd109, 8'd96};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd97};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd132, 8'd120, 8'd106};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd121};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd157, 8'd151, 8'd131};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd136};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd136};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd136};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd161, 8'd155, 8'd131};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd160, 8'd154, 8'd130};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd159, 8'd153, 8'd129};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd159, 8'd153, 8'd130};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd158, 8'd152, 8'd128};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd158, 8'd152, 8'd128};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd158, 8'd152, 8'd130};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd159, 8'd154, 8'd132};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd130};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd130};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd143, 8'd141, 8'd120};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd104};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd92};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd88};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd108, 8'd98, 8'd86};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd108, 8'd98, 8'd86};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd110, 8'd102, 8'd89};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd91};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd93};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd94};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd93};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd90};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd106, 8'd102, 8'd90};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd106, 8'd102, 8'd90};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd103, 8'd90};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd111, 8'd107, 8'd95};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd121, 8'd114, 8'd99};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd129, 8'd121, 8'd106};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd133, 8'd125, 8'd110};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd125, 8'd109};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd110};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd109};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd110};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd112};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd117};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd119};
					endcase
				end
				`ybit'd43: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd83, 8'd99, 8'd70};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd71};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd87, 8'd103, 8'd76};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd73};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd71};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd70};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd70};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd73};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd73};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd86, 8'd99, 8'd73};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd85, 8'd98, 8'd73};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd87, 8'd99, 8'd75};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd90, 8'd103, 8'd74};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd88, 8'd107, 8'd76};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd88, 8'd107, 8'd77};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd87, 8'd103, 8'd76};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd86, 8'd101, 8'd75};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd91, 8'd102, 8'd79};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd91, 8'd103, 8'd81};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd92, 8'd103, 8'd87};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd90, 8'd99, 8'd93};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd88, 8'd99, 8'd103};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd88, 8'd101, 8'd114};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd91, 8'd101, 8'd130};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd92, 8'd102, 8'd137};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd92, 8'd102, 8'd137};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd92, 8'd102, 8'd139};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd93, 8'd101, 8'd139};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd93, 8'd100, 8'd144};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd146};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd151};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd159};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd160};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd162};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd161};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd161};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd160};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd160};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd158};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd156};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd158};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd156};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd152};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd88, 8'd95, 8'd148};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd90, 8'd97, 8'd145};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd90, 8'd97, 8'd146};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd90, 8'd97, 8'd148};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd151};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd156};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd156};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd158};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd158};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd158};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd158};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd157};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd152};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd94, 8'd101, 8'd141};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd95, 8'd102, 8'd129};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd98, 8'd105, 8'd117};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd99, 8'd108, 8'd100};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd102, 8'd108, 8'd88};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd87};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd104, 8'd105, 8'd87};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd104, 8'd106, 8'd85};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd104, 8'd106, 8'd85};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd104, 8'd106, 8'd85};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd85};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd86};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd86};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd110, 8'd103, 8'd87};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd117, 8'd105, 8'd93};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd101};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd116, 8'd112, 8'd108};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd112};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd117};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd117};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd111, 8'd111, 8'd111};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd114, 8'd114, 8'd114};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd115};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd112, 8'd112, 8'd112};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd112, 8'd108, 8'd105};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd114, 8'd105, 8'd100};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd97};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd110, 8'd101, 8'd96};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd110, 8'd100, 8'd91};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd113, 8'd100, 8'd92};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd114, 8'd100, 8'd92};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd113, 8'd100, 8'd91};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd113, 8'd100, 8'd90};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd112, 8'd99, 8'd90};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd114, 8'd101, 8'd92};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd114, 8'd100, 8'd91};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd114, 8'd101, 8'd91};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd113, 8'd101, 8'd91};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd115, 8'd102, 8'd92};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd120, 8'd106, 8'd95};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd125, 8'd109, 8'd96};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd127, 8'd111, 8'd98};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd97};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd124, 8'd108, 8'd95};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd120, 8'd105, 8'd92};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd119, 8'd105, 8'd92};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd119, 8'd105, 8'd92};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd122, 8'd108, 8'd95};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd135, 8'd122, 8'd107};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd123};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd164, 8'd158, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd163, 8'd157, 8'd135};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd163, 8'd157, 8'd136};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd131};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd121};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd125, 8'd124, 8'd103};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd94};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd107, 8'd102, 8'd88};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd86};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd105, 8'd99, 8'd85};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd109, 8'd101, 8'd88};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd89};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd90};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd89};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd88};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd87};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd85};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd84};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd86};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd104, 8'd100, 8'd88};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd114, 8'd104, 8'd92};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd98};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd124, 8'd114, 8'd102};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd123, 8'd118, 8'd106};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd123, 8'd122, 8'd109};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd111};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd112};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd131, 8'd130, 8'd112};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd118};
					endcase
				end
				`ybit'd44: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd69};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd83, 8'd99, 8'd70};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd87, 8'd104, 8'd73};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd89, 8'd106, 8'd76};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd74};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd84, 8'd99, 8'd74};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd73};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd71};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd73};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd86, 8'd99, 8'd73};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd72};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd73};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd87, 8'd97, 8'd76};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd91, 8'd103, 8'd75};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd89, 8'd106, 8'd78};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd85, 8'd104, 8'd76};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd73};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd88, 8'd104, 8'd73};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd91, 8'd104, 8'd75};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd90, 8'd101, 8'd77};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd87, 8'd98, 8'd82};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd86, 8'd97, 8'd89};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd85, 8'd100, 8'd98};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd89, 8'd103, 8'd108};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd90, 8'd104, 8'd112};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd89, 8'd104, 8'd113};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd90, 8'd102, 8'd116};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd89, 8'd101, 8'd115};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd88, 8'd99, 8'd120};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd128};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd142};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd153};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd161};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd160};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd93, 8'd97, 8'd160};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd158};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd157};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd157};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd156};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd156};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd153};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd152};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd88, 8'd95, 8'd144};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd90, 8'd97, 8'd139};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd91, 8'd100, 8'd130};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd92, 8'd100, 8'd130};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd91, 8'd98, 8'd134};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd144};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd151};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd86, 8'd91, 8'd154};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd155};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd157};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd153};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd149};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd142};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd95, 8'd101, 8'd126};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd98, 8'd109, 8'd108};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd100, 8'd108, 8'd89};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd84};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd85};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd102, 8'd104, 8'd83};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd83};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd102, 8'd104, 8'd82};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd84};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd84};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd104, 8'd100, 8'd84};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd87};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd118, 8'd106, 8'd93};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd119, 8'd108, 8'd100};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd114, 8'd109, 8'd106};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd110};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd115};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd115};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd111, 8'd111, 8'd111};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd108};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd100};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd107, 8'd101, 8'd94};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd106, 8'd100, 8'd92};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd109, 8'd99, 8'd93};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd107, 8'd99, 8'd94};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd108, 8'd99, 8'd93};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd107, 8'd97, 8'd91};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd105, 8'd95, 8'd88};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd103, 8'd93, 8'd87};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd103, 8'd93, 8'd87};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd105, 8'd96, 8'd89};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd107, 8'd97, 8'd90};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd106, 8'd96, 8'd90};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd106, 8'd97, 8'd89};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd111, 8'd97, 8'd91};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd117, 8'd103, 8'd91};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd123, 8'd107, 8'd92};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd125, 8'd108, 8'd96};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd126, 8'd109, 8'd97};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd123, 8'd109, 8'd97};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd121, 8'd105, 8'd93};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd114, 8'd102, 8'd91};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd113, 8'd102, 8'd90};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd114, 8'd103, 8'd92};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd124, 8'd111, 8'd99};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd138, 8'd128, 8'd111};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd152, 8'd145, 8'd127};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd134};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd163, 8'd158, 8'd136};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd162, 8'd158, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd161, 8'd158, 8'd135};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd162, 8'd158, 8'd136};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd163, 8'd158, 8'd136};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd128};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd139, 8'd138, 8'd117};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd101};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd94};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd88};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd88};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd85};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd107, 8'd101, 8'd87};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd88};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd88};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd106, 8'd105, 8'd87};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd88};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd87};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd85};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd84};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd85};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd102, 8'd98, 8'd86};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd108, 8'd101, 8'd90};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd113, 8'd105, 8'd92};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd119, 8'd109, 8'd97};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd105};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd109};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd112};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd130, 8'd130, 8'd112};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd135, 8'd133, 8'd116};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd136, 8'd134, 8'd117};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd118};
					endcase
				end
				`ybit'd45: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd68};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd71};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd90, 8'd107, 8'd75};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd93, 8'd110, 8'd74};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd91, 8'd108, 8'd73};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd87, 8'd104, 8'd76};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd83, 8'd102, 8'd73};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd84, 8'd103, 8'd75};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd85, 8'd102, 8'd75};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd89, 8'd99, 8'd74};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd87, 8'd95, 8'd73};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd84, 8'd91, 8'd74};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd85, 8'd94, 8'd75};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd90, 8'd101, 8'd74};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd90, 8'd106, 8'd77};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd85, 8'd104, 8'd76};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd72};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd72};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd71};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd88, 8'd101, 8'd73};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd86, 8'd99, 8'd71};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd84, 8'd96, 8'd74};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd84, 8'd95, 8'd77};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd85};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd91};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd88, 8'd105, 8'd92};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd92};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd91};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd85, 8'd100, 8'd93};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd85, 8'd99, 8'd99};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd87, 8'd96, 8'd109};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd126};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd145};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd158};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd159};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd158};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd158};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd158};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd158};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd156};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd151};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd146};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd88, 8'd96, 8'd134};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd92, 8'd100, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd93, 8'd102, 8'd114};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd93, 8'd102, 8'd114};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd93, 8'd100, 8'd125};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd139};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd86, 8'd91, 8'd148};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd153};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd153};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd154};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd153};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd146};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd93, 8'd100, 8'd131};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd96, 8'd108, 8'd107};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd100, 8'd109, 8'd91};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd100, 8'd105, 8'd83};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd101, 8'd102, 8'd84};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd102, 8'd104, 8'd83};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd84};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd83};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd102, 8'd104, 8'd83};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd101, 8'd102, 8'd84};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd107, 8'd102, 8'd85};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd113, 8'd103, 8'd89};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd119, 8'd107, 8'd93};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd118, 8'd107, 8'd99};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd112, 8'd108, 8'd104};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd109};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd114, 8'd114, 8'd114};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd109, 8'd109, 8'd109};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd105, 8'd101, 8'd97};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd104, 8'd99, 8'd95};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd104, 8'd99, 8'd95};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd96};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd97};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd106, 8'd100, 8'd96};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd103, 8'd97, 8'd93};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd99, 8'd94, 8'd90};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd96, 8'd90, 8'd87};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd96, 8'd91, 8'd87};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd100, 8'd94, 8'd90};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd101, 8'd96, 8'd92};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd101, 8'd96, 8'd92};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd99, 8'd95, 8'd89};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd106, 8'd96, 8'd92};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd113, 8'd100, 8'd91};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd120, 8'd103, 8'd94};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd122, 8'd108, 8'd95};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd123, 8'd109, 8'd96};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd122, 8'd108, 8'd97};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd118, 8'd105, 8'd97};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd112, 8'd103, 8'd95};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd94};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd114, 8'd105, 8'd97};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd124, 8'd116, 8'd104};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd141, 8'd134, 8'd116};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd156, 8'd150, 8'd131};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd135};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd163, 8'd157, 8'd135};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd160, 8'd157, 8'd135};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd161, 8'd158, 8'd136};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd163, 8'd157, 8'd135};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd161, 8'd159, 8'd136};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd131};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd123};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd108};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd97};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd99};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd99, 8'd100, 8'd100};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd100};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd99, 8'd101, 8'd95};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd95};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd96};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd96};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd96};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd99, 8'd100, 8'd97};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd100};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd99};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd95, 8'd96, 8'd98};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd98};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd97};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd101, 8'd97, 8'd97};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd106, 8'd102, 8'd96};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd115, 8'd110, 8'd100};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd107};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd129, 8'd125, 8'd111};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd132, 8'd129, 8'd114};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd136, 8'd133, 8'd116};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd118};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd118};
					endcase
				end
				`ybit'd46: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd70};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd70};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd90, 8'd110, 8'd73};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd94, 8'd115, 8'd74};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd96, 8'd114, 8'd77};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd93, 8'd110, 8'd80};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd89, 8'd108, 8'd76};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd91, 8'd107, 8'd77};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd89, 8'd105, 8'd77};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd90, 8'd99, 8'd74};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd74};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd71};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd87, 8'd90, 8'd72};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd73};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd87, 8'd106, 8'd70};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd86, 8'd105, 8'd73};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd82, 8'd101, 8'd69};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd83, 8'd102, 8'd70};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd82, 8'd101, 8'd72};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd69};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd69};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd69};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd71};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd84, 8'd99, 8'd74};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd75};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd84, 8'd102, 8'd77};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd76};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd84, 8'd99, 8'd75};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd83, 8'd97, 8'd77};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd82, 8'd96, 8'd81};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd82, 8'd94, 8'd94};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd84, 8'd93, 8'd110};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd86, 8'd94, 8'd132};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd153};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd158};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd158};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd158};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd158};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd153};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd141};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd91, 8'd97, 8'd128};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd91, 8'd101, 8'd114};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd92, 8'd104, 8'd105};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd92, 8'd102, 8'd111};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd120};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd136};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd86, 8'd91, 8'd147};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd148};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd91, 8'd98, 8'd131};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd94, 8'd105, 8'd107};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd95, 8'd109, 8'd92};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd99, 8'd106, 8'd83};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd100, 8'd103, 8'd82};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd101, 8'd104, 8'd82};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd102, 8'd106, 8'd83};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd103, 8'd107, 8'd84};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd84};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd83};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd108, 8'd101, 8'd86};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd112, 8'd103, 8'd88};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd117, 8'd105, 8'd91};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd118, 8'd107, 8'd98};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd112, 8'd107, 8'd103};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd109};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd113};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd112, 8'd112, 8'd112};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd109, 8'd109, 8'd109};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd101};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd103, 8'd100, 8'd96};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd104, 8'd100, 8'd96};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd95};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd102};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd102};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd99};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd93};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd89};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd93, 8'd89, 8'd85};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd98, 8'd93, 8'd90};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd94};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd93};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd102, 8'd94, 8'd92};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd102, 8'd96, 8'd87};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd107, 8'd95, 8'd90};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd110, 8'd100, 8'd92};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd117, 8'd107, 8'd98};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd120, 8'd110, 8'd101};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd119, 8'd110, 8'd100};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd116, 8'd105, 8'd99};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd110, 8'd103, 8'd97};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd110, 8'd103, 8'd98};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd104};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd127, 8'd123, 8'd111};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd145, 8'd138, 8'd121};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd158, 8'd152, 8'd127};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd158, 8'd157, 8'd134};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd158, 8'd157, 8'd134};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd128};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd137, 8'd135, 8'd114};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd98};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd106, 8'd107, 8'd97};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd98, 8'd101, 8'd107};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd95, 8'd96, 8'd111};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd114};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd108};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd108};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd96, 8'd101, 8'd108};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd108};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd108};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd111};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd113};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd93, 8'd96, 8'd114};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd92, 8'd94, 8'd112};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd111};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd94, 8'd109};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd96, 8'd98, 8'd105};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd107, 8'd103, 8'd107};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd106};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd109};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd113};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd115};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd118};
					endcase
				end
				`ybit'd47: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd77, 8'd93, 8'd66};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd67};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd73};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd92, 8'd111, 8'd73};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd97, 8'd118, 8'd77};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd99, 8'd117, 8'd74};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd96, 8'd113, 8'd77};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd92, 8'd111, 8'd79};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd91, 8'd107, 8'd78};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd88, 8'd105, 8'd78};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd91, 8'd100, 8'd76};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd86, 8'd94, 8'd76};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd73};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd83, 8'd92, 8'd73};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd84, 8'd99, 8'd71};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd86, 8'd104, 8'd69};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd85, 8'd105, 8'd67};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd83, 8'd102, 8'd69};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd81, 8'd100, 8'd68};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd82, 8'd102, 8'd65};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd67};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd82, 8'd97, 8'd68};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd68};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd66};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd68};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd80, 8'd99, 8'd68};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd81, 8'd100, 8'd69};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd79, 8'd98, 8'd68};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd79, 8'd95, 8'd67};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd78, 8'd95, 8'd68};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd93, 8'd73};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd79, 8'd93, 8'd81};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd82, 8'd93, 8'd99};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd84, 8'd93, 8'd125};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd146};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd153};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd157};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd88, 8'd95, 8'd157};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd157};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd153};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd142};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd91, 8'd97, 8'd133};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd91, 8'd98, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd116};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd88, 8'd96, 8'd120};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd130};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd89, 8'd92, 8'd141};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd147};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd147};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd138};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd91, 8'd101, 8'd114};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd93, 8'd105, 8'd99};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd98, 8'd105, 8'd87};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd96, 8'd104, 8'd81};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd100, 8'd103, 8'd80};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd101, 8'd105, 8'd82};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd101, 8'd105, 8'd82};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd102, 8'd104, 8'd83};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd83};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd107, 8'd99, 8'd83};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd110, 8'd101, 8'd86};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd112, 8'd104, 8'd94};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd111, 8'd105, 8'd100};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd105};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd107};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd112, 8'd112, 8'd112};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd112, 8'd112, 8'd112};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd101};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd104, 8'd100, 8'd100};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd103, 8'd99, 8'd99};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd102};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd103};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd99};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd92};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd88};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd96};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd101};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd99};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd96};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd89};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd100, 8'd92, 8'd90};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd103, 8'd98, 8'd94};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd111, 8'd105, 8'd101};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd116, 8'd111, 8'd107};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd115, 8'd110, 8'd106};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd112, 8'd107, 8'd104};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd104};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd107};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd131, 8'd127, 8'd116};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd149, 8'd143, 8'd125};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd158, 8'd152, 8'd129};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd160, 8'd158, 8'd135};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd159, 8'd157, 8'd134};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd130};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd122};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd128, 8'd126, 8'd105};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd93};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd103, 8'd104, 8'd99};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd97, 8'd98, 8'd110};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd124};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd88, 8'd93, 8'd127};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd123};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd126};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd127};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd127};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd125};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd131};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd132};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd89, 8'd92, 8'd134};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd133};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd131};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd90, 8'd93, 8'd127};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd122};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd112};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd110};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd111};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd113};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd131, 8'd130, 8'd115};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd117};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd117};
					endcase
				end
				`ybit'd48: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd76, 8'd88, 8'd64};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd79, 8'd95, 8'd69};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd84, 8'd102, 8'd70};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd90, 8'd111, 8'd72};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd96, 8'd117, 8'd75};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd97, 8'd118, 8'd74};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd94, 8'd114, 8'd77};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd92, 8'd110, 8'd78};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd91, 8'd107, 8'd77};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd90, 8'd104, 8'd80};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd87, 8'd101, 8'd78};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd85, 8'd97, 8'd78};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd82, 8'd95, 8'd76};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd81, 8'd95, 8'd74};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd72};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd82, 8'd102, 8'd67};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd83, 8'd104, 8'd69};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd82, 8'd102, 8'd63};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd83, 8'd104, 8'd65};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd81, 8'd102, 8'd63};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd80, 8'd100, 8'd63};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd80, 8'd100, 8'd62};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd80, 8'd99, 8'd63};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd64};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd79, 8'd95, 8'd66};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd67};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd67};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd77, 8'd92, 8'd65};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd66};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd79, 8'd92, 8'd66};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd71};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd81};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd94};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd82, 8'd91, 8'd118};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd86, 8'd91, 8'd145};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd154};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd156};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd155};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd156};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd153};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd146};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd86, 8'd93, 8'd139};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd86, 8'd94, 8'd134};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd86, 8'd94, 8'd129};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd86, 8'd93, 8'd135};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd140};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd146};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd154};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd154};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd148};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd141};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd89, 8'd96, 8'd125};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd91, 8'd102, 8'd106};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd97, 8'd104, 8'd91};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd95, 8'd104, 8'd83};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd80};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd80};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd101, 8'd105, 8'd82};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd102, 8'd104, 8'd82};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd100, 8'd102, 8'd81};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd81};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd107, 8'd99, 8'd86};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd106, 8'd102, 8'd90};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd97};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd101};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd90};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd92};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd108};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd107};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd108};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd105};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd106};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd110};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd135, 8'd133, 8'd120};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd149, 8'd147, 8'd126};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd132};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd133};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd131};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd126};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd140, 8'd133, 8'd114};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd98};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd91};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd101, 8'd102, 8'd94};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd97, 8'd100, 8'd109};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd124};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd132};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd134};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd140};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd140};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd84, 8'd91, 8'd138};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd84, 8'd91, 8'd139};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd142};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd142};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd142};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd142};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd138};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd90, 8'd93, 8'd135};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd99, 8'd100, 8'd124};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd118};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd121, 8'd121, 8'd112};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd128, 8'd126, 8'd111};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd131, 8'd130, 8'd112};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd116};
					endcase
				end
				`ybit'd49: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd75, 8'd87, 8'd63};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd68};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd69};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd89, 8'd109, 8'd75};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd95, 8'd115, 8'd78};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd94, 8'd114, 8'd76};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd92, 8'd111, 8'd80};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd90, 8'd108, 8'd82};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd91, 8'd105, 8'd86};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd87};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd85};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd83};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd80};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd97, 8'd78};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd77, 8'd98, 8'd73};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd80, 8'd99, 8'd70};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd80, 8'd102, 8'd67};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd82, 8'd103, 8'd64};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd81, 8'd102, 8'd63};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd81, 8'd102, 8'd63};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd80, 8'd100, 8'd63};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd79, 8'd99, 8'd62};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd77, 8'd97, 8'd61};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd77, 8'd94, 8'd62};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd77, 8'd93, 8'd64};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd75, 8'd91, 8'd64};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd75, 8'd91, 8'd64};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd64};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd76, 8'd88, 8'd64};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd79, 8'd91, 8'd70};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd75};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd86};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd81, 8'd92, 8'd98};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd118};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd144};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd152};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd153};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd155};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd88, 8'd91, 8'd157};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd151};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd148};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd148};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd86, 8'd91, 8'd142};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd148};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd149};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd150};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd152};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd147};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd139};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd89, 8'd97, 8'd121};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd93, 8'd104, 8'd100};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd95, 8'd105, 8'd88};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd97, 8'd101, 8'd78};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd79};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd80};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd99, 8'd101, 8'd79};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd99, 8'd100, 8'd80};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd102, 8'd98, 8'd79};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd83};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd86};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd92};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd98};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd92, 8'd91, 8'd89};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd97};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd108};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd112};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd110};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd105};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd106, 8'd105, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd107};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd113};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd139, 8'd137, 8'd123};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd128};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd153, 8'd151, 8'd131};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd131};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd153, 8'd151, 8'd128};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd119};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd130, 8'd123, 8'd104};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd115, 8'd107, 8'd89};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd111, 8'd102, 8'd85};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd89};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd98, 8'd102, 8'd101};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd96, 8'd102, 8'd113};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd91, 8'd98, 8'd123};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd133};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd140};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd145};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd148};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd150};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd148};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd149};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd143};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd96, 8'd139};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd103, 8'd106, 8'd125};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd118};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd123, 8'd124, 8'd109};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd113};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd110};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd131, 8'd130, 8'd112};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd131, 8'd130, 8'd112};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd132, 8'd131, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
					endcase
				end
				`ybit'd50: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd68};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd80, 8'd95, 8'd73};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd72};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd87, 8'd108, 8'd76};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd90, 8'd111, 8'd78};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd91, 8'd109, 8'd81};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd88, 8'd105, 8'd84};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd91};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd85, 8'd100, 8'd95};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd84, 8'd98, 8'd99};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd83, 8'd97, 8'd100};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd92};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd80, 8'd95, 8'd86};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd79};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd74};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd76, 8'd94, 8'd70};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd78, 8'd97, 8'd66};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd79, 8'd101, 8'd62};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd79, 8'd101, 8'd62};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd80, 8'd102, 8'd63};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd79, 8'd99, 8'd62};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd60};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd77, 8'd94, 8'd59};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd75, 8'd92, 8'd61};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd76, 8'd89, 8'd63};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd61};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd75, 8'd88, 8'd62};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd75, 8'd87, 8'd66};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd77, 8'd88, 8'd70};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd76, 8'd90, 8'd73};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd87};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd100};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd83, 8'd90, 8'd114};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd130};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd144};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd150};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd86, 8'd92, 8'd154};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd153};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd155};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd154};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd150};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd153};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd153};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd153};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd151};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd145};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd129};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd93, 8'd102, 8'd107};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd95, 8'd104, 8'd89};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd93, 8'd102, 8'd77};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd95, 8'd98, 8'd77};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd96, 8'd97, 8'd79};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd97, 8'd99, 8'd78};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd97, 8'd99, 8'd78};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd96, 8'd98, 8'd78};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd97, 8'd98, 8'd80};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd96, 8'd97, 8'd82};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd94, 8'd96, 8'd84};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd93, 8'd94, 8'd88};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd98, 8'd99, 8'd94};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd102};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd102};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd102};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd102};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd110};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd104};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd105};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd123, 8'd123, 8'd112};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd142, 8'd139, 8'd121};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd126};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd153, 8'd151, 8'd128};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd129};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd130};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd157, 8'd155, 8'd132};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd156, 8'd154, 8'd131};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd130};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd130};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd129};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd155, 8'd149, 8'd127};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd148, 8'd145, 8'd124};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd135, 8'd132, 8'd111};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd122, 8'd115, 8'd97};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd112, 8'd100, 8'd86};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd107, 8'd98, 8'd83};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd85};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd103, 8'd104, 8'd93};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd100};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd98, 8'd100, 8'd112};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd123};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd138};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd143};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd148};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd148};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd148};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd148};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd148};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd144};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd138};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd98, 8'd100, 8'd133};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd111, 8'd111, 8'd120};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd122, 8'd118, 8'd110};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd128, 8'd127, 8'd109};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd128, 8'd127, 8'd109};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd110};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd130, 8'd129, 8'd111};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd130, 8'd129, 8'd111};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd130, 8'd129, 8'd111};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd130, 8'd129, 8'd111};
					endcase
				end
				`ybit'd51: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd70};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd83, 8'd98, 8'd75};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd77};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd86, 8'd108, 8'd80};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd87, 8'd107, 8'd85};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd87, 8'd104, 8'd91};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd85, 8'd99, 8'd96};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd82, 8'd96, 8'd106};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd82, 8'd94, 8'd114};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd118};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd81, 8'd92, 8'd116};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd79, 8'd93, 8'd107};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd79, 8'd93, 8'd95};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd92, 8'd85};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd75, 8'd93, 8'd75};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd75, 8'd93, 8'd67};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd76, 8'd95, 8'd62};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd77, 8'd98, 8'd60};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd78, 8'd99, 8'd61};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd78, 8'd99, 8'd61};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd75, 8'd95, 8'd59};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd76, 8'd92, 8'd62};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd74, 8'd89, 8'd60};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd73, 8'd87, 8'd62};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd60};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd74, 8'd86, 8'd59};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd75, 8'd87, 8'd63};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd70};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd78};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd89};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd103};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd119};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd131};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd83, 8'd88, 8'd141};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd150};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd153};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd152};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd153};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd152};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd152};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd153};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd83, 8'd88, 8'd151};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd153};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd151};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd152};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd152};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd148};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd85, 8'd93, 8'd137};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd91, 8'd99, 8'd116};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd91, 8'd104, 8'd94};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd93, 8'd101, 8'd82};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd94, 8'd96, 8'd78};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd77};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd79};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd95, 8'd96, 8'd77};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd77};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd95, 8'd96, 8'd77};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd94, 8'd95, 8'd79};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd79};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd92, 8'd93, 8'd82};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd95, 8'd96, 8'd88};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd99, 8'd101, 8'd94};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd100, 8'd101, 8'd98};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd100, 8'd101, 8'd99};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd102};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd102};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd108};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd105};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd104};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd106};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd128, 8'd128, 8'd113};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd122};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd149, 8'd147, 8'd124};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd127};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd153, 8'd151, 8'd127};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd129};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd130};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd155, 8'd153, 8'd130};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd129};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd154, 8'd152, 8'd129};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd153, 8'd151, 8'd128};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd127};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd152, 8'd149, 8'd126};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd150, 8'd145, 8'd123};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd142, 8'd138, 8'd118};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd128, 8'd124, 8'd104};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd115, 8'd107, 8'd90};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd110, 8'd98, 8'd83};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd107, 8'd96, 8'd82};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd106, 8'd99, 8'd83};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd85};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd89};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd98};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd109};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd86, 8'd89, 8'd130};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd142};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd146};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd146};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd147};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd148};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd147};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd143};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd93, 8'd96, 8'd132};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd106, 8'd107, 8'd125};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd115};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd122, 8'd108};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd126, 8'd126, 8'd108};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd128, 8'd127, 8'd109};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd128, 8'd126, 8'd109};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd108};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd108};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd108};
					endcase
				end
				`ybit'd52: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd77};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd82, 8'd102, 8'd77};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd84, 8'd104, 8'd85};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd84, 8'd104, 8'd93};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd83, 8'd101, 8'd100};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd83, 8'd98, 8'd106};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd115};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd124};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd130};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd135};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd130};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd120};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd79, 8'd91, 8'd104};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd75, 8'd90, 8'd90};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd74, 8'd90, 8'd76};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd67};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd74, 8'd93, 8'd63};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd75, 8'd94, 8'd61};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd76, 8'd96, 8'd63};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd75, 8'd95, 8'd62};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd73, 8'd92, 8'd63};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd63};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd73, 8'd85, 8'd61};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd72, 8'd84, 8'd64};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd61};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd74, 8'd83, 8'd60};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd66};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd75};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd78, 8'd85, 8'd89};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd79, 8'd87, 8'd105};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd119};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd131};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd84, 8'd87, 8'd139};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd144};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd151};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd151};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd153};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd84, 8'd88, 8'd151};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd151};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd83, 8'd88, 8'd150};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd152};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd150};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd152};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd150};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd149};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd82, 8'd89, 8'd142};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd125};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd89, 8'd101, 8'd106};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd91, 8'd102, 8'd91};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd93, 8'd96, 8'd87};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd92, 8'd93, 8'd84};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd92, 8'd94, 8'd85};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd84};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd85};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd92, 8'd98, 8'd83};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd91, 8'd98, 8'd79};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd82};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd82};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd88};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd95, 8'd98, 8'd88};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd97, 8'd100, 8'd90};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd99, 8'd102, 8'd92};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd95};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd99, 8'd100, 8'd93};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd86, 8'd86, 8'd86};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd87, 8'd87, 8'd87};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd102};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd107};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd106};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd102};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd115, 8'd115, 8'd107};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd134, 8'd132, 8'd118};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd123};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd125};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd127};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd125};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd126};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd127};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd127};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd126};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd152, 8'd150, 8'd127};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd125};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd149, 8'd147, 8'd124};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd150, 8'd144, 8'd122};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd119};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd136, 8'd129, 8'd110};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd121, 8'd114, 8'd95};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd101, 8'd84};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd108, 8'd96, 8'd80};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd108, 8'd96, 8'd81};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd108, 8'd96, 8'd82};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd109, 8'd100, 8'd84};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd110, 8'd102, 8'd85};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd105, 8'd101, 8'd89};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd102};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd87, 8'd89, 8'd122};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd136};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd144};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd145};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd146};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd146};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd142};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd137};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd123};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd118};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd124, 8'd121, 8'd110};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd107};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd126, 8'd109};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd125, 8'd124, 8'd106};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd108};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd107};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd105};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd105};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd106};
					endcase
				end
				`ybit'd53: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd83};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd91};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd98};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd107};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd80, 8'd93, 8'd116};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd123};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd130};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd137};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd143};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd144};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd142};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd79, 8'd87, 8'd129};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd113};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd90, 8'd97};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd75, 8'd90, 8'd83};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd73};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd66};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd74, 8'd93, 8'd64};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd74, 8'd93, 8'd66};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd73, 8'd92, 8'd65};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd74, 8'd89, 8'd69};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd72, 8'd86, 8'd69};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd71, 8'd85, 8'd68};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd74, 8'd83, 8'd66};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd63};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd72, 8'd81, 8'd61};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd72, 8'd80, 8'd66};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd81};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd96};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd78, 8'd85, 8'd113};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd124};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd133};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd82, 8'd85, 8'd137};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd82, 8'd85, 8'd140};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd83, 8'd85, 8'd147};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd145};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd150};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd151};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd150};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd151};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd150};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd150};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd148};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd150};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd150};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd150};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd150};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd144};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd82, 8'd91, 8'd132};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd119};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd107};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd100};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd88, 8'd92, 8'd98};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd90, 8'd92, 8'd96};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd93};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd93};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd91, 8'd97, 8'd93};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd90, 8'd97, 8'd92};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd89, 8'd95, 8'd92};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd90, 8'd97, 8'd89};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd92, 8'd97, 8'd83};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd85};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd95, 8'd101, 8'd86};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd95, 8'd102, 8'd87};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd95, 8'd101, 8'd89};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd95, 8'd98, 8'd87};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd88};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd86, 8'd86, 8'd84};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd84, 8'd84, 8'd82};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd92};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd95};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd82};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd84, 8'd84, 8'd84};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd104};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd103};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd103};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd118, 8'd118, 8'd110};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd136, 8'd134, 8'd118};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd122};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd151, 8'd149, 8'd126};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd125};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd150, 8'd148, 8'd120};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd146, 8'd144, 8'd122};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd122};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd124};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd149, 8'd147, 8'd125};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd149, 8'd147, 8'd124};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd149, 8'd143, 8'd122};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd148, 8'd142, 8'd120};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd116};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd137, 8'd132, 8'd112};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd128, 8'd122, 8'd103};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd115, 8'd108, 8'd90};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd98, 8'd82};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd105, 8'd96, 8'd79};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd104, 8'd96, 8'd80};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd108, 8'd94, 8'd81};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd110, 8'd97, 8'd83};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd110, 8'd97, 8'd85};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd106, 8'd97, 8'd88};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd97};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd88, 8'd89, 8'd116};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd131};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd77, 8'd85, 8'd136};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd141};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd145};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd144};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd141};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd129};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd116};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd111};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd124, 8'd123, 8'd106};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd107};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd110};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd108};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd108};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd124, 8'd123, 8'd105};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd104};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd101};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd100};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd101};
					endcase
				end
				`ybit'd54: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd81, 8'd96, 8'd103};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd110};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd80, 8'd92, 8'd116};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd77, 8'd90, 8'd124};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd79, 8'd87, 8'd132};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd135};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd140};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd146};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd138};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd125};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd88, 8'd108};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd76, 8'd89, 8'd96};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd75, 8'd89, 8'd88};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd75, 8'd91, 8'd80};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd74, 8'd90, 8'd78};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd74, 8'd90, 8'd78};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd74, 8'd89, 8'd81};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd83};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd72, 8'd84, 8'd85};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd72, 8'd84, 8'd85};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd79};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd70};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd74, 8'd77, 8'd63};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd74, 8'd75, 8'd69};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd79};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd76, 8'd81, 8'd94};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd78, 8'd86, 8'd106};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd80, 8'd88, 8'd114};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd78, 8'd87, 8'd117};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd125};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd133};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd80, 8'd82, 8'd139};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd143};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd150};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd150};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd149};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd149};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd150};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd149};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd149};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd148};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd148};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd143};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd140};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd82, 8'd89, 8'd132};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd84, 8'd92, 8'd125};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd83, 8'd91, 8'd117};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd118};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd86, 8'd89, 8'd116};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd84, 8'd91, 8'd111};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd111};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd110};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd110};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd86, 8'd94, 8'd109};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd87, 8'd96, 8'd104};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd89, 8'd97, 8'd93};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd92, 8'd100, 8'd89};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd94, 8'd102, 8'd81};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd95, 8'd103, 8'd81};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd94, 8'd100, 8'd84};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd83};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd87, 8'd88, 8'd82};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd83, 8'd84, 8'd78};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd84, 8'd85, 8'd78};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd85, 8'd86, 8'd81};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd90, 8'd91, 8'd86};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd92, 8'd93, 8'd88};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd83, 8'd83, 8'd83};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd80, 8'd80, 8'd80};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd82};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd101};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd100};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd119, 8'd118, 8'd110};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd118};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd122};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd149, 8'd147, 8'd124};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd124};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd120};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd140, 8'd137, 8'd119};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd116};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd141, 8'd138, 8'd120};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd121};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd120};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd143, 8'd137, 8'd115};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd139, 8'd133, 8'd111};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd137, 8'd126, 8'd106};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd131, 8'd122, 8'd103};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd122, 8'd110, 8'd94};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd114, 8'd102, 8'd86};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd109, 8'd97, 8'd81};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd105, 8'd96, 8'd79};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd103, 8'd97, 8'd80};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd107, 8'd92, 8'd79};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd108, 8'd94, 8'd81};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd108, 8'd95, 8'd83};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd103, 8'd96, 8'd82};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd92};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd105};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd115};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd125};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd131};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd137};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd80, 8'd82, 8'd140};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd86, 8'd89, 8'd135};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd121};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd109};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd105};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd122, 8'd122, 8'd104};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd107};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd126, 8'd125, 8'd107};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd110};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd132, 8'd129, 8'd112};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd132, 8'd130, 8'd112};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd127, 8'd126, 8'd108};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd124, 8'd121, 8'd106};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd101};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd99};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd98};
					endcase
				end
				`ybit'd55: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd117};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd123};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd77, 8'd86, 8'd130};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd137};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd139};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd144};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd146};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd149};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd150};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd149};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd142};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd131};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd86, 8'd118};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd111};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd76, 8'd87, 8'd102};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd76, 8'd88, 8'd99};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd76, 8'd89, 8'd98};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd75, 8'd88, 8'd97};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd96};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd99};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd75, 8'd83, 8'd102};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd74, 8'd82, 8'd101};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd91};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd76};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd74, 8'd76, 8'd68};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd73, 8'd76, 8'd67};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd74, 8'd76, 8'd73};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd84};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd76, 8'd87, 8'd92};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd94};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd102};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd78, 8'd85, 8'd112};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd127};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd139};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd144};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd148};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd141};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd140};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd135};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd135};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd132};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd130};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd129};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd129};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd129};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd129};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd81, 8'd89, 8'd126};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd82, 8'd91, 8'd120};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd85, 8'd96, 8'd106};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd91, 8'd95, 8'd98};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd92};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd89, 8'd98, 8'd92};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd88};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd86, 8'd93, 8'd85};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd82};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd77};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd77};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd82};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd82};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd84};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd91, 8'd93, 8'd91};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd80, 8'd80, 8'd80};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd78, 8'd78, 8'd78};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd97};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd109};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd137, 8'd135, 8'd119};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd145, 8'd143, 8'd119};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd148, 8'd146, 8'd124};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd144, 8'd142, 8'd121};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd118};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd126, 8'd128, 8'd112};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd113};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd114};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd120};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd115};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd136, 8'd128, 8'd108};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd128, 8'd120, 8'd101};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd125, 8'd115, 8'd96};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd121, 8'd109, 8'd93};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd118, 8'd103, 8'd88};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd116, 8'd99, 8'd85};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd97, 8'd81};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd106, 8'd96, 8'd80};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd102, 8'd93, 8'd77};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd101, 8'd91, 8'd77};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd103, 8'd91, 8'd79};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd100, 8'd89, 8'd77};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd97, 8'd93, 8'd81};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd93, 8'd96, 8'd82};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd90, 8'd95, 8'd91};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd84, 8'd93, 8'd101};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd83, 8'd91, 8'd110};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd121};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd129};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd134};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd126};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd98, 8'd100, 8'd114};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd110, 8'd106, 8'd104};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd97};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd100};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd124, 8'd121, 8'd104};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd125, 8'd124, 8'd106};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd110};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd134, 8'd131, 8'd112};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd136, 8'd133, 8'd114};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd133, 8'd130, 8'd111};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd129, 8'd126, 8'd108};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd101};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd118, 8'd114, 8'd97};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd96};
					endcase
				end
				`ybit'd56: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd131};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd136};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd142};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd145};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd146};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd149};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd149};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd149};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd143};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd140};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd134};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd128};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd123};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd77, 8'd85, 8'd121};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd119};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd118};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd74, 8'd83, 8'd117};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd119};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd116};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd115};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd102};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd82};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd75, 8'd78, 8'd70};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd75, 8'd78, 8'd69};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd76, 8'd79, 8'd71};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd73};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd76, 8'd90, 8'd77};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd91, 8'd78};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd87};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd106};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd125};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd138};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd144};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd146};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd146};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd146};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd144};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd143};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd142};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd142};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd140};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd142};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd141};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd140};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd140};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd139};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd140};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd133};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd123};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd83, 8'd90, 8'd115};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd109};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd83, 8'd88, 8'd107};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd82, 8'd89, 8'd105};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd100};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd89};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd84, 8'd92, 8'd83};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd88, 8'd91, 8'd76};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd86, 8'd94, 8'd74};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd88, 8'd95, 8'd78};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd88, 8'd95, 8'd79};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd88, 8'd91, 8'd83};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd87, 8'd87, 8'd87};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd83, 8'd83, 8'd83};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd79};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd78, 8'd78, 8'd78};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd96};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd98};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd104};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd122, 8'd122, 8'd112};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd119};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd143, 8'd140, 8'd121};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd141, 8'd138, 8'd121};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd128, 8'd126, 8'd113};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd109};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd112};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd134, 8'd132, 8'd118};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd141, 8'd138, 8'd118};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd138, 8'd131, 8'd113};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd127, 8'd119, 8'd103};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd118, 8'd108, 8'd94};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd119, 8'd102, 8'd90};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd116, 8'd99, 8'd85};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd114, 8'd98, 8'd83};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd112, 8'd96, 8'd81};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd109, 8'd97, 8'd81};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd106, 8'd95, 8'd79};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd102, 8'd92, 8'd78};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd99, 8'd90, 8'd76};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd94, 8'd87, 8'd73};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd93, 8'd88, 8'd73};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd94, 8'd91, 8'd73};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd75};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd90, 8'd96, 8'd82};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd85};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd87, 8'd92, 8'd95};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd105};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd117};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd84, 8'd85, 8'd121};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd90, 8'd91, 8'd115};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd101};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd94};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd95};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd115, 8'd112, 8'd96};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd100};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd124, 8'd124, 8'd106};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd108};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd134, 8'd131, 8'd112};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd138, 8'd135, 8'd116};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd115};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd132, 8'd129, 8'd113};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd125, 8'd122, 8'd105};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd99};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd95};
					endcase
				end
				`ybit'd57: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd139};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd142};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd145};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd80, 8'd84, 8'd147};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd148};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd140};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd139};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd136};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd133};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd131};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd131};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd77, 8'd80, 8'd129};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd128};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd122};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd110};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd95};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd80};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd68};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd64};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd78, 8'd86, 8'd67};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd70};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd68};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd74};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd77, 8'd91, 8'd86};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd106};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd127};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd141};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd144};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd144};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd80, 8'd82, 8'd139};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd80, 8'd82, 8'd139};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd141};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd144};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd145};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd79, 8'd80, 8'd144};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd78, 8'd79, 8'd143};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd76, 8'd81, 8'd137};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd132};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd129};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd128};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd126};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd120};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd114};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd81, 8'd86, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd92};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd81};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd88, 8'd97, 8'd74};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd73};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd77};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd80};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd86, 8'd87, 8'd82};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd86, 8'd86, 8'd86};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd89};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd84, 8'd84, 8'd84};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd76, 8'd76, 8'd76};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd76, 8'd76, 8'd76};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd82};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd95};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd96};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd104};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd125, 8'd125, 8'd113};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd137, 8'd137, 8'd118};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd117};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd116};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd112};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd110};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd110};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd113};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd132, 8'd132, 8'd118};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd137, 8'd136, 8'd118};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd109};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd120, 8'd112, 8'd100};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd114, 8'd100, 8'd91};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd113, 8'd98, 8'd86};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd114, 8'd96, 8'd84};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd112, 8'd94, 8'd81};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd113, 8'd94, 8'd81};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd111, 8'd95, 8'd80};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd109, 8'd95, 8'd78};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd101, 8'd93, 8'd75};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd94, 8'd91, 8'd72};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd71};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd71};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd91, 8'd93, 8'd71};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd74};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd91, 8'd94, 8'd73};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd88, 8'd96, 8'd80};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd84};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd85, 8'd91, 8'd96};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd109};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd110};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd92, 8'd93, 8'd103};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd96};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd89};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd90};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd95};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd103};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd125, 8'd122, 8'd105};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd127, 8'd124, 8'd107};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd131, 8'd128, 8'd108};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd135, 8'd132, 8'd113};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd115};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd133, 8'd130, 8'd111};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd124, 8'd123, 8'd105};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd97};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd93};
					endcase
				end
				`ybit'd58: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd143};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd145};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd146};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd147};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd146};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd142};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd138};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd136};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd77, 8'd80, 8'd130};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd76, 8'd81, 8'd121};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd110};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd77, 8'd86, 8'd98};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd85};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd77, 8'd86, 8'd74};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd75, 8'd88, 8'd67};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd77, 8'd91, 8'd65};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd78, 8'd92, 8'd67};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd77, 8'd94, 8'd67};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd70};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd79, 8'd95, 8'd76};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd76, 8'd90, 8'd91};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd112};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd132};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd144};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd143};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd143};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd139};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd140};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd140};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd138};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd134};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd128};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd127};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd131};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd138};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd139};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd139};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd140};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd143};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd144};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd145};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd77, 8'd78, 8'd143};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd76, 8'd78, 8'd142};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd145};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd140};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd140};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd75, 8'd78, 8'd136};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd77, 8'd79, 8'd136};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd75, 8'd78, 8'd133};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd128};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd119};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd80, 8'd88, 8'd106};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd89};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd89, 8'd99, 8'd77};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd88, 8'd99, 8'd70};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd72};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd83, 8'd90, 8'd74};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd84, 8'd86, 8'd76};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd84, 8'd86, 8'd79};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd87, 8'd88, 8'd83};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd88};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd82};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd77, 8'd77, 8'd77};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd74};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd76, 8'd76, 8'd76};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd97};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd110, 8'd110, 8'd105};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd125, 8'd125, 8'd112};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd114};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd128, 8'd127, 8'd113};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd111};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd107};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd107};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd107};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd112};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd117};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd107};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd111, 8'd107, 8'd98};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd109, 8'd99, 8'd92};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd110, 8'd94, 8'd82};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd112, 8'd95, 8'd83};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd112, 8'd94, 8'd80};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd112, 8'd94, 8'd80};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd111, 8'd95, 8'd80};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd108, 8'd94, 8'd78};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd103, 8'd94, 8'd77};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd74};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd94, 8'd90, 8'd71};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd72};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd91, 8'd92, 8'd72};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd90, 8'd92, 8'd71};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd89, 8'd92, 8'd71};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd89, 8'd92, 8'd72};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd87, 8'd90, 8'd74};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd86, 8'd88, 8'd84};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd87, 8'd88, 8'd98};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd90, 8'd91, 8'd101};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd96};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd88};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd94, 8'd93, 8'd86};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd89};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd95};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd101};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd103};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd106};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd127, 8'd124, 8'd106};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd129, 8'd126, 8'd107};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd131, 8'd128, 8'd109};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd106};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd119, 8'd118, 8'd100};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd88};
					endcase
				end
				`ybit'd59: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd77, 8'd80, 8'd144};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd144};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd144};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd144};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd145};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd138};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd136};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd131};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd123};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd113};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd100};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd79, 8'd91, 8'd86};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd77, 8'd92, 8'd75};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd77, 8'd92, 8'd72};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd77, 8'd93, 8'd66};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd79, 8'd95, 8'd68};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd69};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd71};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd76};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd78, 8'd92, 8'd90};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd75, 8'd86, 8'd105};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd122};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd135};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd82, 8'd137};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd139};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd135};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd133};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd134};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd132};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd78, 8'd85, 8'd131};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd129};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd129};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd124};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd119};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd112};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd112};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd119};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd79, 8'd87, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd125};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd130};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd132};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd139};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd143};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd144};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd144};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd142};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd141};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd142};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd142};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd140};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd138};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd134};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd129};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd117};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd99};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd83};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd88, 8'd97, 8'd76};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd85, 8'd94, 8'd74};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd75};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd84, 8'd87, 8'd75};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd83, 8'd85, 8'd75};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd85, 8'd86, 8'd78};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd86, 8'd87, 8'd81};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd84, 8'd85, 8'd79};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd78};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd78, 8'd78, 8'd76};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd74};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd71, 8'd71, 8'd71};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd74};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd92};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd90};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd91};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd93, 8'd93, 8'd93};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd94};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd107};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd109};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd116, 8'd116, 8'd106};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd104};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd102};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd103};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd109, 8'd110, 8'd105};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd111};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd113};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd110};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd104};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd99};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd107, 8'd97, 8'd94};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd108, 8'd94, 8'd83};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd108, 8'd94, 8'd81};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd110, 8'd92, 8'd79};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd110, 8'd92, 8'd78};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd92, 8'd78};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd110, 8'd94, 8'd79};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd106, 8'd92, 8'd76};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd99, 8'd93, 8'd75};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd99, 8'd91, 8'd74};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd97, 8'd91, 8'd74};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd93, 8'd89, 8'd73};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd70};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd69};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd70};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd84, 8'd86, 8'd72};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd85, 8'd87, 8'd78};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd87, 8'd91, 8'd89};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd94};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd89};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd87};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd87};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd93};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd98};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd103};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd103};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd123, 8'd122, 8'd104};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd123, 8'd122, 8'd104};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd103};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd101};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd98};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd92};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd85};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd82};
					endcase
				end
				`ybit'd60: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd140};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd76, 8'd81, 8'd143};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd136};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd132};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd127};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd112};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd99};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd79, 8'd94, 8'd87};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd75};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd78, 8'd96, 8'd71};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd66};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd66};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd66};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd71};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd77, 8'd96, 8'd76};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd76, 8'd92, 8'd91};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd74, 8'd86, 8'd104};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd72, 8'd81, 8'd118};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd70, 8'd78, 8'd131};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd134};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd134};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd126};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd75, 8'd83, 8'd124};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd123};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd123};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd119};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd115};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd81, 8'd90, 8'd112};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd81, 8'd90, 8'd111};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd106};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd99};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd93};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd93};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd80, 8'd92, 8'd98};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd105};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd80, 8'd88, 8'd110};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd79, 8'd87, 8'd115};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd124};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd134};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd140};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd140};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd141};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd139};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd139};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd139};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd141};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd141};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd136};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd125};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd107};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd95};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd84, 8'd90, 8'd85};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd83, 8'd90, 8'd81};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd80};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd85, 8'd88, 8'd74};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd71};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd72};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd73};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd72};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd77, 8'd78, 8'd73};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd73, 8'd74, 8'd71};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd70, 8'd71, 8'd69};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd68, 8'd68, 8'd67};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd73, 8'd73, 8'd74};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd80};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd87, 8'd87, 8'd87};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd87, 8'd87, 8'd87};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd88};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd87, 8'd87, 8'd87};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd90};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd95, 8'd94, 8'd93};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd96};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd100};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd103};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd106, 8'd105, 8'd100};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd102};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd99};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd98};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd100};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd106};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd106};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd103};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd101};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd97};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd102, 8'd94, 8'd93};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd103, 8'd92, 8'd85};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd106, 8'd90, 8'd80};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd108, 8'd89, 8'd77};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd107, 8'd89, 8'd77};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd108, 8'd89, 8'd77};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd106, 8'd90, 8'd75};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd106, 8'd90, 8'd76};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd104, 8'd90, 8'd75};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd101, 8'd89, 8'd73};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd98, 8'd87, 8'd74};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd93, 8'd83, 8'd73};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd88, 8'd79, 8'd69};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd85, 8'd78, 8'd67};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd82, 8'd78, 8'd65};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd68};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd88, 8'd85, 8'd74};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd83};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd87};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd92, 8'd91, 8'd85};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd85};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd88};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd96};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd99};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd102};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd101};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd101};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd101};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd99};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd93};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd86};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd80};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd76};
					endcase
				end
				`ybit'd61: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd143};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd136};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd128};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd116};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd78, 8'd91, 8'd100};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd80, 8'd95, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd81, 8'd98, 8'd79};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd74};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd79, 8'd99, 8'd73};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd73};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd78, 8'd97, 8'd75};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd75};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd77, 8'd93, 8'd82};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd75, 8'd90, 8'd93};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd73, 8'd86, 8'd104};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd71, 8'd80, 8'd119};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd69, 8'd77, 8'd126};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd70, 8'd77, 8'd132};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd133};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd82, 8'd120};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd111};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd106};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd77, 8'd90, 8'd101};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd100};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd80, 8'd91, 8'd97};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd80, 8'd94, 8'd94};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd82, 8'd95, 8'd91};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd84, 8'd96, 8'd92};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd84, 8'd97, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd84, 8'd98, 8'd84};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd83, 8'd98, 8'd76};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd83, 8'd98, 8'd76};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd83};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd83, 8'd96, 8'd85};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd90};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd80, 8'd91, 8'd95};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd78, 8'd85, 8'd112};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd125};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd137};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd138};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd143};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd137};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd138};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd139};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd140};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd141};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd140};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd129};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd119};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd110};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd106};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd78, 8'd85, 8'd101};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd81, 8'd87, 8'd93};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd84};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd80};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd76};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd79, 8'd82, 8'd74};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd73};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd74, 8'd76, 8'd71};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd72, 8'd74, 8'd69};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd69, 8'd72, 8'd65};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd69, 8'd70, 8'd64};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd69};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd77, 8'd79, 8'd74};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd82};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd84, 8'd84, 8'd84};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd85, 8'd85, 8'd85};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd87, 8'd87, 8'd87};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd90, 8'd90, 8'd88};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd94, 8'd95, 8'd89};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd94};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd96};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd96};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd96};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd98, 8'd99, 8'd95};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd97, 8'd98, 8'd93};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd96};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd96};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd98};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd99};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd96};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd94};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd92};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd100, 8'd92, 8'd90};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd99, 8'd90, 8'd83};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd101, 8'd89, 8'd78};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd102, 8'd87, 8'd75};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd101, 8'd87, 8'd74};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd101, 8'd87, 8'd74};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd104, 8'd88, 8'd73};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd104, 8'd88, 8'd74};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd102, 8'd87, 8'd74};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd98, 8'd84, 8'd73};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd94, 8'd82, 8'd70};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd89, 8'd78, 8'd68};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd85, 8'd75, 8'd65};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd80, 8'd71, 8'd64};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd82, 8'd73, 8'd66};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd84, 8'd79, 8'd68};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd91, 8'd86, 8'd74};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd82};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd92, 8'd91, 8'd86};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd91, 8'd91, 8'd83};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd87};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd93};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd98};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd101};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd101};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd100};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd100};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd99};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd96};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd89};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd83};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd77};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd73};
					endcase
				end
				`ybit'd62: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd142};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd140};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd70, 8'd77, 8'd139};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd134};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd127};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd76, 8'd89, 8'd109};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd80, 8'd95, 8'd94};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd84};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd79, 8'd98, 8'd80};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd78, 8'd96, 8'd84};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd76, 8'd94, 8'd83};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd75, 8'd93, 8'd81};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd76, 8'd94, 8'd82};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd75, 8'd92, 8'd87};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd75, 8'd89, 8'd98};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd72, 8'd83, 8'd105};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd118};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd69, 8'd77, 8'd124};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd129};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd71, 8'd76, 8'd131};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd126};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd75, 8'd84, 8'd109};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd93};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd79, 8'd92, 8'd86};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd80, 8'd94, 8'd82};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd81, 8'd94, 8'd82};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd83};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd82, 8'd96, 8'd77};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd84, 8'd100, 8'd74};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd74};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd73};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd85, 8'd102, 8'd70};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd81, 8'd100, 8'd69};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd69};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd69};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd83, 8'd99, 8'd72};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd84, 8'd96, 8'd73};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd81, 8'd92, 8'd78};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd78, 8'd86, 8'd100};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd116};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd134};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd140};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd142};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd138};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd137};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd136};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd137};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd141};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd140};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd134};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd130};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd121};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd74, 8'd77, 8'd121};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd115};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd110};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd100};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd91};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd82};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd80};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd73, 8'd76, 8'd78};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd73, 8'd74, 8'd77};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd71, 8'd73, 8'd69};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd64};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd67};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd72, 8'd75, 8'd68};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd76, 8'd79, 8'd72};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd79, 8'd80, 8'd76};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd79, 8'd80, 8'd76};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd80, 8'd81, 8'd77};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd80, 8'd81, 8'd77};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd81, 8'd82, 8'd78};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd79};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd84, 8'd84, 8'd81};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd85};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd94, 8'd96, 8'd89};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd91};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd95};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd96};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd107, 8'd107, 8'd96};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd97};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd95};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd94};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd95};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd96};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd97};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd97};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd95};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd92};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd90};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd95, 8'd94, 8'd89};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd100, 8'd93, 8'd85};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd98, 8'd90, 8'd79};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd100, 8'd88, 8'd76};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd101, 8'd88, 8'd76};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd102, 8'd87, 8'd76};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd102, 8'd87, 8'd76};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd101, 8'd87, 8'd76};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd100, 8'd85, 8'd74};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd97, 8'd82, 8'd71};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd91, 8'd78, 8'd70};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd85, 8'd74, 8'd66};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd79, 8'd69, 8'd60};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd76, 8'd67, 8'd62};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd78, 8'd70, 8'd64};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd84, 8'd80, 8'd68};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd90, 8'd86, 8'd74};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd80};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd89, 8'd88, 8'd83};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd84};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd99, 8'd100, 8'd86};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd92};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd117, 8'd116, 8'd98};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd99};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd99};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd99};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd99};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd116, 8'd116, 8'd98};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd96};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd91};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd87};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd81};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd80};
					endcase
				end
				`ybit'd63: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd140};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd72, 8'd75, 8'd139};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd140};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd140};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd135};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd73, 8'd82, 8'd122};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd76, 8'd89, 8'd104};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd78, 8'd94, 8'd90};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd78, 8'd95, 8'd89};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd74, 8'd89, 8'd95};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd73, 8'd87, 8'd101};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd72, 8'd85, 8'd104};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd72, 8'd85, 8'd104};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd72, 8'd85, 8'd103};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd72, 8'd84, 8'd108};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd115};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd70, 8'd77, 8'd118};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd69, 8'd77, 8'd125};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd69, 8'd78, 8'd119};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd118};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd117};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd111};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd76, 8'd89, 8'd94};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd80, 8'd91, 8'd76};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd79, 8'd95, 8'd70};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd68};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd68};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd78, 8'd98, 8'd67};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd66};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd65};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd66};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd66};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd83, 8'd101, 8'd64};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd82, 8'd102, 8'd64};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd82, 8'd102, 8'd64};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd64};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd67};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd84, 8'd97, 8'd69};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd74};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd75, 8'd86, 8'd93};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd71, 8'd80, 8'd114};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd71, 8'd76, 8'd133};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd138};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd136};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd137};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd136};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd136};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd137};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd71, 8'd76, 8'd140};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd139};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd139};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd134};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd71, 8'd76, 8'd133};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd134};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd134};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd69, 8'd76, 8'd128};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd70, 8'd78, 8'd124};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd116};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd108};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd100};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd98};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd93};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd90};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd84};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd75};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd75, 8'd78, 8'd68};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd77, 8'd80, 8'd72};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd76, 8'd78, 8'd71};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd77, 8'd78, 8'd69};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd78, 8'd79, 8'd70};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd79, 8'd80, 8'd71};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd79, 8'd80, 8'd71};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd78, 8'd79, 8'd71};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd81, 8'd82, 8'd76};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd86, 8'd87, 8'd80};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd94, 8'd95, 8'd88};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd92};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd99};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd105};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd106};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd125, 8'd120, 8'd106};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd123, 8'd119, 8'd102};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd105};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd115, 8'd116, 8'd103};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd104};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd104};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd102};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd106, 8'd105, 8'd101};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd100};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd99};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd96};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd95};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd102, 8'd96, 8'd88};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd99, 8'd96, 8'd83};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd100, 8'd92, 8'd79};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd101, 8'd93, 8'd80};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd102, 8'd93, 8'd80};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd102, 8'd93, 8'd80};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd101, 8'd92, 8'd80};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd99, 8'd89, 8'd77};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd96, 8'd87, 8'd74};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd90, 8'd83, 8'd72};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd85, 8'd75, 8'd66};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd79, 8'd68, 8'd60};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd76, 8'd67, 8'd62};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd78, 8'd69, 8'd64};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd85, 8'd79, 8'd72};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd89, 8'd85, 8'd77};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd82};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd88, 8'd87, 8'd82};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd88};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd105, 8'd106, 8'd91};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd96};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd117, 8'd116, 8'd98};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd118, 8'd115, 8'd98};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd97};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd97};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd97};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd97};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd97};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd93};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd89};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd85};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd83};
					endcase
				end
				`ybit'd64: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd138};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd137};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd136};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd124};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd73, 8'd85, 8'd106};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd75, 8'd88, 8'd100};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd72, 8'd86, 8'd99};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd70, 8'd81, 8'd111};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd115};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd117};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd119};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd119};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd120};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd69, 8'd76, 8'd122};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd69, 8'd76, 8'd120};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd70, 8'd78, 8'd116};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd107};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd73, 8'd84, 8'd103};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd101};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd96};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd78, 8'd91, 8'd83};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd80, 8'd95, 8'd72};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd79, 8'd98, 8'd66};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd65};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd81, 8'd98, 8'd65};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd64};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd60};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd81, 8'd98, 8'd62};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd81, 8'd98, 8'd62};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd64};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd64};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd83, 8'd97, 8'd63};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd77};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd96};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd69, 8'd77, 8'd115};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd131};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd133};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd136};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd135};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd135};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd137};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd135};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd131};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd127};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd69, 8'd76, 8'd120};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd117};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd68, 8'd71, 8'd111};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd67, 8'd70, 8'd109};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd66, 8'd69, 8'd104};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd99};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd86};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd80};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd74};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd75, 8'd79, 8'd75};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd73};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd78, 8'd80, 8'd72};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd79, 8'd82, 8'd69};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd65};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd80, 8'd83, 8'd67};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd85, 8'd87, 8'd72};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd93, 8'd96, 8'd81};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd92};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd103};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd110};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd132, 8'd130, 8'd113};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd115};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd135, 8'd135, 8'd111};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd136, 8'd135, 8'd116};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd135, 8'd134, 8'd115};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd116};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd118};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd113, 8'd113, 8'd116};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd108, 8'd110, 8'd116};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd107, 8'd109, 8'd114};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd109, 8'd109, 8'd111};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd108, 8'd108, 8'd111};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd106, 8'd105, 8'd110};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd103};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd98};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd103, 8'd100, 8'd92};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd103, 8'd98, 8'd89};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd106, 8'd100, 8'd92};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd105, 8'd99, 8'd90};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd105, 8'd99, 8'd91};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd106, 8'd98, 8'd89};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd106, 8'd97, 8'd89};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd102, 8'd94, 8'd85};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd97, 8'd88, 8'd81};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd90, 8'd81, 8'd74};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd83, 8'd74, 8'd66};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd75, 8'd70, 8'd64};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd75, 8'd72, 8'd67};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd72};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd75};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd77};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd88, 8'd87, 8'd83};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd88};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd92};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd96};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd97};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd94};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd94};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd91};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd90};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd90};
					endcase
				end
				`ybit'd65: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd138};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd138};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd134};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd125};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd71, 8'd79, 8'd118};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd69, 8'd80, 8'd110};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd67, 8'd76, 8'd115};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd73, 8'd121};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd65, 8'd72, 8'd126};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd130};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd131};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd132};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd66, 8'd73, 8'd131};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd128};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd69, 8'd76, 8'd118};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd71, 8'd82, 8'd102};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd74, 8'd88, 8'd93};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd76, 8'd91, 8'd84};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd83};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd79, 8'd92, 8'd81};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd77, 8'd93, 8'd68};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd78, 8'd95, 8'd60};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd77, 8'd97, 8'd60};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd81, 8'd98, 8'd61};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd61};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd65};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd60};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd62};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd62};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd60};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd83, 8'd101, 8'd63};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd64};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd65};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd83, 8'd96, 8'd68};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd81};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd72, 8'd80, 8'd102};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd119};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd131};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd131};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd136};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd134};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd134};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd137};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd136};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd130};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd129};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd64, 8'd70, 8'd125};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd120};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd120};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd64, 8'd71, 8'd115};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd68, 8'd75, 8'd103};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd96};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd93};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd91};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd86};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd78};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd69};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd66};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd85, 8'd88, 8'd66};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd71};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd83};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd98};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd129, 8'd128, 8'd108};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd115};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd134, 8'd132, 8'd119};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd135, 8'd133, 8'd121};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd137, 8'd134, 8'd124};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd138, 8'd136, 8'd123};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd139, 8'd137, 8'd124};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd133, 8'd130, 8'd124};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd128};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd107, 8'd110, 8'd129};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd129};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd128};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd128};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd103, 8'd104, 8'd128};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd101, 8'd103, 8'd124};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd100, 8'd103, 8'd118};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd113};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd101, 8'd101, 8'd105};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd104};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd103};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd103};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd101};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd100};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd105, 8'd101, 8'd99};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd104, 8'd100, 8'd98};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd92};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd96, 8'd92, 8'd88};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd88, 8'd84, 8'd80};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd81, 8'd76, 8'd70};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd77, 8'd74, 8'd69};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd76, 8'd75, 8'd72};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd76};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd80};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd84};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd90};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd94};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd95};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd89};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd90};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd90};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd91};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd94};
					endcase
				end
				`ybit'd66: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd136};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd137};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd130};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd124};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd123};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd125};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd127};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd134};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd134};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd135};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd125};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd69, 8'd78, 8'd111};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd74, 8'd85, 8'd92};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd77, 8'd91, 8'd80};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd77, 8'd94, 8'd73};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd72};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd75, 8'd93, 8'd69};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd76, 8'd95, 8'd64};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd76, 8'd95, 8'd63};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd77, 8'd98, 8'd59};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd79, 8'd100, 8'd61};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd80, 8'd100, 8'd61};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd61};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd82, 8'd99, 8'd62};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd64};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd87, 8'd101, 8'd65};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd86, 8'd100, 8'd65};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd80, 8'd96, 8'd69};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd75, 8'd86, 8'd86};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd70, 8'd77, 8'd106};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd121};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd132};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd135};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd135};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd136};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd127};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd125};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd124};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd117};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd114};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd110};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd108};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd101};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd92};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd81};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd74};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd68};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd74};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd101, 8'd107, 8'd86};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd121, 8'd121, 8'd101};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd130, 8'd130, 8'd116};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd118};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd121, 8'd121, 8'd122};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd119, 8'd119, 8'd126};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd121, 8'd120, 8'd129};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd124, 8'd124, 8'd127};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd124, 8'd125, 8'd128};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd130};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd107, 8'd109, 8'd132};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd95, 8'd99, 8'd134};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd136};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd87, 8'd93, 8'd134};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd88, 8'd95, 8'd134};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd89, 8'd92, 8'd131};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd88, 8'd93, 8'd125};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd88, 8'd91, 8'd119};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd90, 8'd91, 8'd115};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd90, 8'd92, 8'd112};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd91, 8'd93, 8'd113};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd92, 8'd93, 8'd111};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd111};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd95, 8'd94, 8'd110};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd96, 8'd96, 8'd105};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd105};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd98, 8'd97, 8'd103};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd98};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd88};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd88, 8'd84, 8'd80};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd77, 8'd77, 8'd71};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd73, 8'd72, 8'd70};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd75, 8'd74, 8'd73};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd80, 8'd80, 8'd80};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd87, 8'd88, 8'd82};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd86};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd90};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd91};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd91};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd90};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd90};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd89};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd88};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd88};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd89};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd91};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd94};
					endcase
				end
				`ybit'd67: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd135};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd135};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd135};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd135};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd137};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd135};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd132};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd66, 8'd69, 8'd134};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd134};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd135};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd133};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd123};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd70, 8'd79, 8'd109};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd85};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd77, 8'd93, 8'd71};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd77, 8'd96, 8'd64};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd77, 8'd97, 8'd60};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd76, 8'd95, 8'd63};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd73, 8'd93, 8'd58};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd74, 8'd93, 8'd59};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd78, 8'd98, 8'd60};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd78, 8'd99, 8'd60};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd80, 8'd101, 8'd62};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd61};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd83, 8'd100, 8'd62};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd84, 8'd101, 8'd63};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd86, 8'd101, 8'd64};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd84, 8'd98, 8'd63};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd80, 8'd95, 8'd69};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd75, 8'd86, 8'd86};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd68, 8'd76, 8'd107};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd122};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd134};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd134};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd135};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd133};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd134};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd68, 8'd71, 8'd134};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd68, 8'd71, 8'd133};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd132};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd131};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd133};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd133};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd133};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd133};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd131};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd130};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd128};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd65, 8'd68, 8'd126};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd124};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd124};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd63, 8'd70, 8'd117};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd106};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd93};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd89};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd82, 8'd85, 8'd86};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd86, 8'd88, 8'd85};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd93};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd112, 8'd112, 8'd108};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd122, 8'd122, 8'd118};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd124};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd127};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd98, 8'd99, 8'd130};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd98, 8'd101, 8'd132};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd98, 8'd103, 8'd133};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd101, 8'd104, 8'd132};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd99, 8'd102, 8'd132};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd137};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd83, 8'd89, 8'd139};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd77, 8'd85, 8'd143};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd142};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd142};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd140};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd138};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd134};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd131};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd79, 8'd82, 8'd127};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd124};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd121};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd79, 8'd83, 8'd120};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd80, 8'd83, 8'd117};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd82, 8'd85, 8'd115};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd87, 8'd89, 8'd111};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd91, 8'd93, 8'd108};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd109};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd102};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd95};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd90, 8'd89, 8'd84};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd74};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd73, 8'd73, 8'd71};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd75, 8'd74, 8'd73};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd79};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd84, 8'd85, 8'd81};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd86};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd88};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd91};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd92};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd92};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd93};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd113, 8'd112, 8'd93};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd92};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd90};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd87};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd84};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd84};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd86};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd87};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd90};
					endcase
				end
				`ybit'd68: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd134};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd134};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd134};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd65, 8'd72, 8'd134};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd134};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd134};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd133};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd133};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd133};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd122};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd108};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd73, 8'd88, 8'd82};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd76, 8'd94, 8'd67};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd77, 8'd97, 8'd60};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd77, 8'd98, 8'd59};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd75, 8'd95, 8'd58};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd75, 8'd95, 8'd58};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd75, 8'd95, 8'd58};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd75, 8'd95, 8'd58};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd78, 8'd99, 8'd60};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd80, 8'd101, 8'd62};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd83, 8'd101, 8'd61};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd62};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd78, 8'd96, 8'd58};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd84, 8'd98, 8'd63};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd84, 8'd98, 8'd63};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd69};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd72};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd78, 8'd91, 8'd75};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd73, 8'd84, 8'd88};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd67, 8'd76, 8'd106};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd64, 8'd71, 8'd121};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd69, 8'd71, 8'd129};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd69, 8'd70, 8'd129};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd69, 8'd72, 8'd123};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd121};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd123};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd126};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd131};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd129};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd127};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd126};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd122};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd124};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd124};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd126};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd126};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd126};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd129};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd125};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd125};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd123};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd66, 8'd69, 8'd118};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd107};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd71, 8'd76, 8'd101};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd98};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd76, 8'd78, 8'd100};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd82, 8'd85, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd113};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd103, 8'd106, 8'd122};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd128};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd88, 8'd94, 8'd128};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd134};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd134};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd134};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd82, 8'd89, 8'd138};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd137};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd137};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd138};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd139};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd139};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd72, 8'd81, 8'd138};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd139};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd138};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd135};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd132};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd129};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd126};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd122};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd80, 8'd82, 8'd119};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd112};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd87, 8'd86, 8'd108};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd92, 8'd94, 8'd106};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd103};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd101};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd92};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd91, 8'd90, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd73};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd74};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd76, 8'd76, 8'd76};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd78, 8'd78, 8'd78};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd79};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd82};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd94, 8'd93, 8'd84};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd87};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd89};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd91};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd94};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd95};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd116, 8'd115, 8'd95};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd114, 8'd111, 8'd94};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd90};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd86};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd83};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd83};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd83};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd84};
					endcase
				end
				`ybit'd69: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd133};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd66, 8'd71, 8'd133};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd133};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd132};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd132};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd133};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd132};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd131};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd132};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd128};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd119};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd71, 8'd80, 8'd103};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd78};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd75, 8'd92, 8'd64};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd76, 8'd94, 8'd58};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd58};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd75, 8'd94, 8'd57};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd94, 8'd57};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd73, 8'd93, 8'd56};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd77, 8'd94, 8'd58};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd78, 8'd96, 8'd58};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd61};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd60};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd81, 8'd97, 8'd62};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd79, 8'd94, 8'd69};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd78, 8'd91, 8'd77};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd73, 8'd88, 8'd81};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd71, 8'd85, 8'd85};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd69, 8'd80, 8'd95};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd65, 8'd73, 8'd112};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd125};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd131};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd67, 8'd69, 8'd132};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd66, 8'd69, 8'd132};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd122};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd110};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd73, 8'd77, 8'd108};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd112};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd123};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd67, 8'd68, 8'd133};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd131};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd129};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd128};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd128};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd128};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd128};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd128};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd61, 8'd64, 8'd127};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd123};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd122};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd63, 8'd66, 8'd121};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd117};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd115};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd115};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd71, 8'd73, 8'd113};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd117};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd118};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd120};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd120};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd120};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd120};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd65, 8'd72, 8'd118};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd67, 8'd71, 8'd115};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd115};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd69, 8'd73, 8'd114};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd110};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd111};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd112};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd118};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd127};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd129};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd130};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd135};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd139};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd136};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd138};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd137};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd139};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd143};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd142};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd143};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd142};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd138};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd132};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd128};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd87, 8'd90, 8'd124};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd90, 8'd94, 8'd122};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd94, 8'd95, 8'd117};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd112};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd105};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd102};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd96};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd98, 8'd98, 8'd88};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd89, 8'd88, 8'd81};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd73};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd75, 8'd75, 8'd73};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd76, 8'd76, 8'd75};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd77, 8'd77, 8'd77};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd77};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd79};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd80};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd99, 8'd96, 8'd84};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd86};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd88};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd93};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd97};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd99};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd98};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd94};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd90};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd86};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd82};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd96, 8'd94, 8'd79};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd79};
					endcase
				end
				`ybit'd70: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd132};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd131};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd126};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd66, 8'd74, 8'd114};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd94};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd72};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd74, 8'd90, 8'd59};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd72, 8'd91, 8'd54};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd72, 8'd92, 8'd55};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd72, 8'd92, 8'd55};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd75, 8'd92, 8'd56};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd56};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd78, 8'd96, 8'd58};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd63};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd78, 8'd93, 8'd67};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd74, 8'd87, 8'd75};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd90};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd98};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd101};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd66, 8'd73, 8'd111};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd119};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd128};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd132};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd67, 8'd68, 8'd132};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd133};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd128};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd113};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd101};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd93};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd101};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd118};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd66, 8'd68, 8'd128};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd127};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd124};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd117};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd62, 8'd69, 8'd114};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd63, 8'd72, 8'd110};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd107};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd67, 8'd75, 8'd99};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd72, 8'd80, 8'd96};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd76, 8'd81, 8'd93};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd93};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd96};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd77, 8'd80, 8'd97};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd98};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd99};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd76, 8'd78, 8'd102};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd75, 8'd78, 8'd103};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd102};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd106};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd108};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd70, 8'd77, 8'd108};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd108};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd108};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd111};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd114};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd76, 8'd81, 8'd119};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd121};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd123};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd127};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd130};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd135};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd137};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd137};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd138};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd143};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd72, 8'd80, 8'd142};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd141};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd138};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd132};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd80, 8'd88, 8'd129};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd97, 8'd100, 8'd124};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd108, 8'd110, 8'd122};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd118};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd111};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd107};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd120, 8'd115, 8'd104};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd114, 8'd110, 8'd97};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd103, 8'd100, 8'd87};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd88, 8'd88, 8'd81};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd72};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd78, 8'd78, 8'd76};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd79};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd79};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd77};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd78};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd86, 8'd86, 8'd77};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd83};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd85};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd87};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd92};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd94};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd98};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd100};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd100};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd117, 8'd116, 8'd96};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd91};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd85};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd78};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd77};
					endcase
				end
				`ybit'd71: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd128};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd131};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd131};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd131};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd125};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd66, 8'd74, 8'd110};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd70, 8'd81, 8'd87};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd68};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd72, 8'd88, 8'd58};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd72, 8'd88, 8'd56};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd73, 8'd90, 8'd55};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd71, 8'd91, 8'd54};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd71, 8'd91, 8'd54};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd73, 8'd90, 8'd54};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd76, 8'd93, 8'd57};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd57};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd80, 8'd98, 8'd60};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd80, 8'd97, 8'd62};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd80, 8'd93, 8'd64};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd72, 8'd89, 8'd71};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd67, 8'd80, 8'd88};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd62, 8'd70, 8'd102};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd59, 8'd67, 8'd109};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd114};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd60, 8'd67, 8'd119};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd126};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd132};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd124};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd111};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd71, 8'd79, 8'd94};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd85};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd69, 8'd77, 8'd96};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd65, 8'd72, 8'd116};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd126};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd59, 8'd62, 8'd126};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd121};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd111};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd66, 8'd73, 8'd100};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd68, 8'd76, 8'd92};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd90};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd82};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd79};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd77};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd82, 8'd89, 8'd77};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd79};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd80};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd83};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd82, 8'd86, 8'd83};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd80, 8'd86, 8'd85};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd82, 8'd88, 8'd87};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd82, 8'd87, 8'd88};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd81, 8'd85, 8'd88};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd93};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd94};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd92};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd77, 8'd80, 8'd96};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd75, 8'd83, 8'd99};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd103};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd75, 8'd83, 8'd100};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd76, 8'd84, 8'd103};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd74, 8'd85, 8'd107};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd114};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd123};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd130};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd136};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd74, 8'd79, 8'd142};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd143};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd70, 8'd78, 8'd140};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd138};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd67, 8'd78, 8'd133};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd78, 8'd84, 8'd126};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd96, 8'd100, 8'd120};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd117, 8'd117, 8'd123};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd120};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd117};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd111};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd128, 8'd125, 8'd107};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd98};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd105, 8'd101, 8'd89};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd78};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd81, 8'd80, 8'd77};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd79};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd87, 8'd86, 8'd82};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd88, 8'd87, 8'd83};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd85, 8'd84, 8'd79};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd79};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd81};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd79};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd83};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd85};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd87};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd89};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd115, 8'd112, 8'd93};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd97};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd100};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd101};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd97};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd94};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd101, 8'd97, 8'd85};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd79};
					endcase
				end
				`ybit'd72: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd117};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd118};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd119};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd124};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd124};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd124};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd124};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd125};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd62, 8'd65, 8'd128};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd130};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd60, 8'd67, 8'd128};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd60, 8'd67, 8'd129};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd124};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd64, 8'd72, 8'd109};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd90};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd69, 8'd81, 8'd74};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd70, 8'd84, 8'd65};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd65};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd72, 8'd88, 8'd59};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd70, 8'd91, 8'd53};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd71, 8'd91, 8'd54};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd72, 8'd89, 8'd53};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd73, 8'd90, 8'd54};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd73, 8'd90, 8'd54};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd76, 8'd94, 8'd56};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd78, 8'd96, 8'd58};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd59};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd79, 8'd96, 8'd58};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd78, 8'd95, 8'd64};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd77, 8'd89, 8'd70};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd68, 8'd81, 8'd82};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd62, 8'd71, 8'd98};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd115};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd121};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd122};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd127};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd130};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd131};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd127};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd118};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd66, 8'd73, 8'd99};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd68, 8'd76, 8'd94};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd66, 8'd73, 8'd102};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd118};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd62, 8'd65, 8'd129};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd62, 8'd65, 8'd129};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd130};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd127};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd117};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd107};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd85};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd76};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd72};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd68};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd66};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd84, 8'd95, 8'd62};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd85, 8'd96, 8'd65};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd84, 8'd95, 8'd66};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd84, 8'd95, 8'd66};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd83, 8'd92, 8'd67};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd83, 8'd91, 8'd69};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd68};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd69};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd71};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd85, 8'd94, 8'd72};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd85, 8'd94, 8'd74};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd84, 8'd93, 8'd73};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd82, 8'd91, 8'd75};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd76};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd77};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd80};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd79, 8'd85, 8'd81};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd83};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd83};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd80, 8'd89, 8'd91};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd103};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd77, 8'd85, 8'd117};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd132};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd136};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd142};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd141};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd69, 8'd78, 8'd140};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd135};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd126};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd89, 8'd91, 8'd122};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd111, 8'd110, 8'd122};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd130, 8'd128, 8'd117};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd119};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd142, 8'd135, 8'd114};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd134, 8'd132, 8'd108};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd100};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd90};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd80};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd86, 8'd86, 8'd76};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd91, 8'd92, 8'd82};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd87};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd97, 8'd97, 8'd87};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd92, 8'd92, 8'd81};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd79};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd79};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd78};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd81};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd103, 8'd99, 8'd83};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd84};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd105, 8'd101, 8'd88};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd85};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd89};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd95};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd100};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd101};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd118, 8'd115, 8'd96};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd110, 8'd106, 8'd88};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd100, 8'd100, 8'd80};
					endcase
				end
				`ybit'd73: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd99};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd99};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd105};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd62, 8'd69, 8'd112};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd116};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd116};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd119};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd121};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd60, 8'd65, 8'd122};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd62, 8'd67, 8'd124};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd114};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd63, 8'd74, 8'd98};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd65, 8'd78, 8'd88};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd79};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd67, 8'd83, 8'd73};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd69, 8'd86, 8'd65};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd73, 8'd89, 8'd59};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd54};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd73, 8'd90, 8'd54};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd74, 8'd88, 8'd54};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd76, 8'd90, 8'd55};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd77, 8'd91, 8'd57};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd76, 8'd93, 8'd59};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd75, 8'd93, 8'd61};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd75, 8'd91, 8'd66};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd73, 8'd88, 8'd68};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd70, 8'd83, 8'd75};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd63, 8'd74, 8'd93};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd59, 8'd66, 8'd110};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd119};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd126};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd127};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd129};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd130};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd126};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd119};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd62, 8'd70, 8'd110};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd106};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd111};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd120};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd126};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd130};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd128};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd117};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd100};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd79};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd80, 8'd89, 8'd68};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd80, 8'd89, 8'd63};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd60};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd83, 8'd92, 8'd62};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd61};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd60};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd60};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd60};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd61};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd85, 8'd94, 8'd61};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd62};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd89, 8'd98, 8'd65};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd89, 8'd99, 8'd65};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd64};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd89, 8'd98, 8'd65};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd64};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd83, 8'd94, 8'd65};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd85, 8'd93, 8'd66};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd83, 8'd91, 8'd64};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd81, 8'd89, 8'd67};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd79, 8'd86, 8'd65};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd80, 8'd87, 8'd68};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd81, 8'd90, 8'd71};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd83, 8'd92, 8'd74};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd85, 8'd92, 8'd87};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd103};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd74, 8'd83, 8'd126};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd136};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd136};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd140};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd136};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd137};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd137};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd71, 8'd80, 8'd137};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd137};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd136};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd136};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd136};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd67, 8'd74, 8'd128};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd123};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd94, 8'd95, 8'd121};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd117, 8'd116, 8'd117};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd115};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd139, 8'd137, 8'd115};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd137, 8'd130, 8'd111};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd99};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd88};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd95, 8'd94, 8'd82};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd84};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd89};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd95};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd94};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd89};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd84};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd96, 8'd94, 8'd80};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd82};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd99, 8'd96, 8'd79};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd81};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd82};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd83};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd83};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd84};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd89};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd93};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd98};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd98};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd96};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd91};
					endcase
				end
				`ybit'd74: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd59, 8'd72, 8'd77};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd60, 8'd74, 8'd78};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd59, 8'd71, 8'd83};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd95};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd101};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd62, 8'd70, 8'd104};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd60, 8'd67, 8'd106};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd59, 8'd66, 8'd110};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd117};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd126};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd61, 8'd64, 8'd128};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd123};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd60, 8'd66, 8'd117};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd61, 8'd68, 8'd112};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd62, 8'd70, 8'd104};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd96};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd64, 8'd78, 8'd83};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd68, 8'd85, 8'd69};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd72, 8'd88, 8'd60};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd55};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd77, 8'd91, 8'd56};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd77, 8'd91, 8'd56};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd76, 8'd90, 8'd62};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd72, 8'd87, 8'd65};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd70, 8'd84, 8'd71};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd69, 8'd82, 8'd75};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd68, 8'd79, 8'd79};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd64, 8'd73, 8'd91};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd59, 8'd67, 8'd104};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd119};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd122};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd124};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd126};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd127};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd60, 8'd66, 8'd128};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd62, 8'd65, 8'd129};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd62, 8'd65, 8'd129};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd62, 8'd65, 8'd129};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd129};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd124};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd123};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd122};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd118};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd124};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd61, 8'd63, 8'd129};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd61, 8'd67, 8'd129};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd127};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd125};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd123};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd113};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd65, 8'd72, 8'd96};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd74};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd60};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd55};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd55};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd57};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd60};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd84, 8'd95, 8'd54};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd85, 8'd96, 8'd55};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd85, 8'd96, 8'd55};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd87, 8'd97, 8'd60};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd61};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd88, 8'd98, 8'd61};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd87, 8'd97, 8'd59};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd86, 8'd97, 8'd59};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd83, 8'd95, 8'd56};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd81, 8'd90, 8'd58};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd55};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd58};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd57};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd82, 8'd93, 8'd60};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd71};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd88};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd112};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd131};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd135};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd139};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd136};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd137};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd70, 8'd79, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd137};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd72, 8'd79, 8'd137};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd70, 8'd77, 8'd135};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd138};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd64, 8'd72, 8'd129};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd68, 8'd74, 8'd127};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd124};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd97, 8'd99, 8'd117};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd116};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd130, 8'd127, 8'd111};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd132, 8'd126, 8'd107};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd98};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd89};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd89};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd97};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd123, 8'd122, 8'd102};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd102};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd122, 8'd118, 8'd99};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd91};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd86};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd85};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd86};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd85};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd81};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd81};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd79};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd79};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd82};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd87};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd111, 8'd108, 8'd90};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd95};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd98};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd94};
					endcase
				end
				`ybit'd75: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd59, 8'd73, 8'd57};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd59, 8'd73, 8'd57};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd62};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd75};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd60, 8'd73, 8'd85};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd60, 8'd71, 8'd87};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd91};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd96};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd57, 8'd64, 8'd105};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd116};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd121};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd126};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd122};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd116};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd115};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd106};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd64, 8'd75, 8'd91};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd67, 8'd82, 8'd75};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd71, 8'd87, 8'd62};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd74, 8'd90, 8'd58};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd59};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd74, 8'd91, 8'd57};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd75, 8'd92, 8'd57};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd75, 8'd91, 8'd63};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd67};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd65, 8'd80, 8'd75};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd61, 8'd74, 8'd87};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd61, 8'd72, 8'd92};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd98};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd59, 8'd66, 8'd105};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd115};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd120};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd124};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd62, 8'd66, 8'd129};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd128};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd128};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd60, 8'd66, 8'd128};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd126};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd125};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd60, 8'd66, 8'd128};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd127};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd125};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd123};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd115};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd64, 8'd71, 8'd94};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd66};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd57};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd55};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd56};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd59};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd57};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd86, 8'd96, 8'd59};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd86, 8'd97, 8'd57};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd58};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd58};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd56};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd58};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd58};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd56};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd54};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd54};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd57};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd85, 8'd95, 8'd67};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd83, 8'd92, 8'd83};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd77, 8'd83, 8'd106};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd126};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd67, 8'd72, 8'd131};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd137};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd70, 8'd76, 8'd137};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd133};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd135};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd132};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd133};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd133};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd131};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd72, 8'd78, 8'd130};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd127};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd125};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd72, 8'd76, 8'd125};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd121};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd116};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd109};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd121, 8'd117, 8'd102};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd96};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd87};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd114, 8'd112, 8'd95};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd127, 8'd125, 8'd102};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd135, 8'd132, 8'd108};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd138, 8'd132, 8'd108};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd135, 8'd129, 8'd107};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd130, 8'd124, 8'd101};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd125, 8'd120, 8'd97};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd97};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd118, 8'd115, 8'd96};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd114, 8'd111, 8'd92};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd88};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd83};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd80};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd77};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd77};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd96, 8'd94, 8'd79};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd82};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd87};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd114, 8'd113, 8'd92};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd95};
					endcase
				end
				`ybit'd76: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd44};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd41};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd56, 8'd68, 8'd46};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd59};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd58, 8'd70, 8'd73};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd76};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd76};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd80};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd90};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd104};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd115};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd121};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd124};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd125};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd126};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd60, 8'd63, 8'd126};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd126};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd123};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd123};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd120};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd59, 8'd66, 8'd112};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd98};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd66, 8'd79, 8'd82};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd68, 8'd83, 8'd74};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd68, 8'd84, 8'd67};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd69, 8'd85, 8'd65};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd70, 8'd85, 8'd63};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd64};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd69, 8'd84, 8'd69};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd65, 8'd78, 8'd76};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd60, 8'd71, 8'd89};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd109};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd111};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd115};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd122};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd122};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd127};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd125};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd127};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd127};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd125};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd125};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd126};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd126};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd125};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd126};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd122};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd121};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd121};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd122};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd122};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd113};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd89};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd65};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd56};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd54};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd77, 8'd85, 8'd54};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd80, 8'd88, 8'd54};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd57};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd56};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd86, 8'd95, 8'd58};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd84, 8'd95, 8'd57};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd57};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd56};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd55};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd52};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd52};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd53};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd82, 8'd91, 8'd56};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd82, 8'd93, 8'd64};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd80, 8'd89, 8'd79};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd71, 8'd82, 8'd103};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd64, 8'd73, 8'd120};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd128};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd131};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd133};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd67, 8'd73, 8'd135};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd73, 8'd78, 8'd131};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd130};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd86, 8'd90, 8'd125};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd88, 8'd91, 8'd123};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd85, 8'd89, 8'd124};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd123};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd84, 8'd86, 8'd124};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd81, 8'd84, 8'd123};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd79, 8'd82, 8'd122};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd76, 8'd80, 8'd120};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd117};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd91, 8'd96, 8'd113};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd106, 8'd105, 8'd106};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd97};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd92};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd88};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd89};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd94};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd131, 8'd127, 8'd102};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd112};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd112};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd144, 8'd139, 8'd111};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd142, 8'd137, 8'd109};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd140, 8'd134, 8'd107};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd136, 8'd132, 8'd107};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd107};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd129, 8'd124, 8'd103};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd122, 8'd117, 8'd96};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd91};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd85};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd78};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd73};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd74};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd75};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd76};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd81};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd87};
					endcase
				end
				`ybit'd77: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd55, 8'd69, 8'd36};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd40};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd53, 8'd67, 8'd52};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd54, 8'd66, 8'd61};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd54, 8'd66, 8'd61};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd59};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd64};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd72};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd83};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd97};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd111};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd119};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd124};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd120};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd117};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd60, 8'd65, 8'd118};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd117};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd60, 8'd66, 8'd118};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd118};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd118};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd118};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd119};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd118};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd57, 8'd64, 8'd111};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd100};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd63, 8'd75, 8'd89};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd64, 8'd77, 8'd81};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd63, 8'd78, 8'd75};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd64, 8'd78, 8'd76};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd66, 8'd77, 8'd78};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd66, 8'd77, 8'd79};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd64, 8'd75, 8'd84};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd91};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd101};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd52, 8'd59, 8'd111};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd117};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd119};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd119};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd121};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd123};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd57, 8'd64, 8'd126};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd57, 8'd64, 8'd126};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd124};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd125};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd127};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd125};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd125};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd59, 8'd63, 8'd126};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd125};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd124};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd123};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd124};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd121};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd121};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd53, 8'd61, 8'd107};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd59, 8'd66, 8'd84};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd62};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd72, 8'd81, 8'd53};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd52};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd52};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd77, 8'd84, 8'd50};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd55};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd54};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd54};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd54};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd84, 8'd94, 8'd57};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd54};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd54};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd53};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd52};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd52};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd56};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd63};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd79, 8'd88, 8'd79};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd66, 8'd79, 8'd101};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd116};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd121};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd58, 8'd67, 8'd126};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd62, 8'd69, 8'd127};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd65, 8'd72, 8'd130};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd72, 8'd77, 8'd126};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd84, 8'd87, 8'd124};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd96, 8'd98, 8'd118};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd98, 8'd101, 8'd113};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd95, 8'd98, 8'd112};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd94, 8'd95, 8'd112};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd95, 8'd97, 8'd113};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd98, 8'd100, 8'd116};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd95, 8'd97, 8'd115};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd91, 8'd93, 8'd113};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd90, 8'd92, 8'd112};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd95, 8'd98, 8'd106};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd102};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd99};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd114, 8'd111, 8'd92};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd89};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd90};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd97};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd132, 8'd127, 8'd103};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd113};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd150, 8'd145, 8'd116};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd149, 8'd144, 8'd115};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd147, 8'd141, 8'd117};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd145, 8'd139, 8'd112};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd141, 8'd135, 8'd110};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd133, 8'd127, 8'd104};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd95};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd89};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd81};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd74};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd71};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd70};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd71};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd75};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd96, 8'd94, 8'd79};
					endcase
				end
				`ybit'd78: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd34};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd36};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd51, 8'd63, 8'd41};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd46};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd51};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd49};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd48};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd52};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd58};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd67};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd53, 8'd60, 8'd80};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd101};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd113};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd120};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd56, 8'd59, 8'd124};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd118};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd124};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd55, 8'd58, 8'd124};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd121};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd118};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd61, 8'd64, 8'd114};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd108};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd104};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd106};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd108};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd61, 8'd66, 8'd109};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd60, 8'd65, 8'd108};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd114};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd113};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd110};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd109};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd97};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd60, 8'd71, 8'd90};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd63, 8'd72, 8'd83};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd82};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd62, 8'd71, 8'd82};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd59, 8'd71, 8'd88};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd93};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd97};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd102};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd112};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd54, 8'd57, 8'd121};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd123};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd58, 8'd61, 8'd124};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd125};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd57, 8'd60, 8'd123};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd124};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd122};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd121};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd117};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd105};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd80};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd67, 8'd70, 8'd57};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd51};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd71, 8'd75, 8'd52};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd51};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd49};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd52};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd54};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd55};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd55};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd53};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd56};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd82, 8'd92, 8'd55};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd53};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd53};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd50};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd54};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd81, 8'd91, 8'd64};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd77};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd68, 8'd79, 8'd96};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd63, 8'd70, 8'd114};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd59, 8'd67, 8'd123};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd123};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd66, 8'd72, 8'd125};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd127};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd77, 8'd81, 8'd125};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd85, 8'd90, 8'd115};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd110};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd102};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd103, 8'd99, 8'd98};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd95};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd100};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd110, 8'd109, 8'd106};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd107};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd103};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd102, 8'd102, 8'd106};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd106, 8'd106, 8'd104};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd117, 8'd114, 8'd106};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd123, 8'd120, 8'd103};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd127, 8'd122, 8'd99};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd126, 8'd120, 8'd98};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd97};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd97};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd136, 8'd130, 8'd106};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd145, 8'd139, 8'd115};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd150, 8'd145, 8'd116};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd150, 8'd145, 8'd116};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd149, 8'd144, 8'd115};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd149, 8'd144, 8'd115};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd149, 8'd144, 8'd114};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd113};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd140, 8'd135, 8'd111};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd129, 8'd127, 8'd102};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd97};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd88};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd75};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd89, 8'd85, 8'd72};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd67};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd64};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd67};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd72};
					endcase
				end
				`ybit'd79: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd53, 8'd67, 8'd33};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd35};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd40};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd44};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd45};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd39};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd51, 8'd63, 8'd38};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd42};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd45};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd49};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd62};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd84};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd53, 8'd60, 8'd102};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd114};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd55, 8'd58, 8'd119};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd117};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd119};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd57, 8'd60, 8'd121};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd117};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd112};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd62, 8'd68, 8'd100};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd74, 8'd88};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd64, 8'd75, 8'd82};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd63, 8'd76, 8'd82};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd63, 8'd75, 8'd85};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd64, 8'd72, 8'd90};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd63, 8'd72, 8'd90};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd95};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd98};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd98};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd97};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd59, 8'd71, 8'd88};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd60, 8'd72, 8'd83};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd61, 8'd73, 8'd74};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd61, 8'd73, 8'd73};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd79};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd88};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd100};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd104};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd109};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd113};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd115};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd116};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd118};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd57, 8'd61, 8'd124};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd120};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd118};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd118};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd118};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd51, 8'd57, 8'd116};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd100};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd57, 8'd63, 8'd75};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd51};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd48};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd49};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd65, 8'd70, 8'd47};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd69, 8'd76, 8'd46};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd49};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd53};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd53};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd80, 8'd90, 8'd53};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd52};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd50};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd53};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd57};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd69};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd71, 8'd83, 8'd88};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd66, 8'd75, 8'd105};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd70, 8'd75, 8'd115};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd115};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd117};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd83, 8'd87, 8'd119};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd87, 8'd89, 8'd114};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd110};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd103, 8'd99, 8'd100};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd90};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd89};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd105, 8'd100, 8'd88};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd91};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd114, 8'd110, 8'd95};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd114, 8'd110, 8'd94};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd93};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd92};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd93};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd100};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd131, 8'd129, 8'd106};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd137, 8'd133, 8'd104};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd137, 8'd131, 8'd103};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd134, 8'd133, 8'd103};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd135, 8'd133, 8'd108};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd141, 8'd136, 8'd111};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd147, 8'd141, 8'd117};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd150, 8'd145, 8'd116};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd149, 8'd144, 8'd115};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd115};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd112};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd134, 8'd132, 8'd107};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd125, 8'd124, 8'd98};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd96};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd83};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd94, 8'd90, 8'd77};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd68};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd61};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd62};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd66};
					endcase
				end
				`ybit'd80: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd34};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd39};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd41};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd37};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd36};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd38};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd38};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd40};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd40};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd52};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd50, 8'd58, 8'd71};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd92};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd104};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd111};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd115};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd114};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd114};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd109};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd62, 8'd69, 8'd98};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd86};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd80, 8'd72};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd65, 8'd81, 8'd67};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd65, 8'd81, 8'd66};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd67, 8'd80, 8'd68};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd67, 8'd80, 8'd71};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd67, 8'd79, 8'd76};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd66, 8'd78, 8'd78};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd67, 8'd78, 8'd79};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd66, 8'd77, 8'd80};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd65, 8'd76, 8'd80};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd63, 8'd75, 8'd75};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd63, 8'd75, 8'd71};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd63, 8'd74, 8'd63};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd63};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd64, 8'd73, 8'd69};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd61, 8'd72, 8'd79};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd89};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd93};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd99};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd103};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd106};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd113};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd119};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd119};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd123};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd122};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd120};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd117};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd118};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd119};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd118};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd112};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd97};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd61, 8'd61, 8'd73};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd65, 8'd68, 8'd55};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd68, 8'd72, 8'd47};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd66, 8'd69, 8'd48};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd66, 8'd67, 8'd46};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd65, 8'd71, 8'd49};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd48};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd49};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd50};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd49};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd53};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd53};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd53};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd54};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd63};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd76};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd95};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd78, 8'd83, 8'd112};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd114};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd116};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd113};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd103, 8'd103, 8'd109};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd105};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd103, 8'd100, 8'd95};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd88};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd83};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd84};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd88};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd112, 8'd111, 8'd90};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd88};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd84};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd100, 8'd98, 8'd82};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd88};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd116, 8'd113, 8'd93};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd132, 8'd125, 8'd104};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd140, 8'd134, 8'd110};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd112};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd112};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd142, 8'd135, 8'd112};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd116};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd149, 8'd143, 8'd119};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd149, 8'd143, 8'd119};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd112};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd111};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd143, 8'd139, 8'd109};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd139, 8'd133, 8'd109};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd132, 8'd126, 8'd102};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd125, 8'd118, 8'd98};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd114, 8'd108, 8'd88};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd79};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd87, 8'd86, 8'd69};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd64};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd61};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd66};
					endcase
				end
				`ybit'd81: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd47, 8'd61, 8'd31};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd33};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd37};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd33};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd37};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd35};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd37};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd36};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd38};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd38};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd49};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd61};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd77};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd88};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd97};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd101};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd57, 8'd65, 8'd103};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd58, 8'd67, 8'd100};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd94};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd63, 8'd74, 8'd79};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd68, 8'd81, 8'd69};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd66, 8'd84, 8'd57};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd66, 8'd86, 8'd52};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd85, 8'd52};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd68, 8'd85, 8'd54};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd69, 8'd86, 8'd52};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd69, 8'd85, 8'd58};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd69, 8'd85, 8'd61};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd69, 8'd85, 8'd61};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd68, 8'd83, 8'd62};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd67, 8'd82, 8'd60};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd65, 8'd81, 8'd56};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd64, 8'd79, 8'd56};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd65, 8'd78, 8'd52};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd66, 8'd79, 8'd53};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd66, 8'd78, 8'd58};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd64, 8'd78, 8'd60};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd63, 8'd75, 8'd71};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd62, 8'd74, 8'd78};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd82};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd64, 8'd69, 8'd87};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd91};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd107};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd115};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd54, 8'd57, 8'd121};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd117};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd116};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd116};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd117};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd116};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd115};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd118};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd106};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd93};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd59, 8'd61, 8'd66};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd63, 8'd67, 8'd49};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd66, 8'd70, 8'd45};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd68, 8'd65, 8'd45};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd63, 8'd63, 8'd43};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd63, 8'd69, 8'd47};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd71, 8'd77, 8'd46};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd48};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd49};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd50};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd50};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd52};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd53};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd80, 8'd92, 8'd54};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd78, 8'd90, 8'd67};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd74, 8'd83, 8'd84};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd83, 8'd86, 8'd99};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd98, 8'd100, 8'd105};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd111};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd118, 8'd117, 8'd109};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd114, 8'd114, 8'd102};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd112, 8'd108, 8'd96};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd90};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd81};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd85};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd89};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd92};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd93};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd88};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd81};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd78};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd80};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd84};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd123, 8'd117, 8'd95};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd132, 8'd126, 8'd102};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd135, 8'd129, 8'd106};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd136, 8'd130, 8'd106};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd137, 8'd131, 8'd106};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd141, 8'd135, 8'd111};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd145, 8'd139, 8'd115};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd116};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd112};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd111};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd110};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd139, 8'd133, 8'd109};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd135, 8'd129, 8'd105};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd128, 8'd121, 8'd101};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd121, 8'd114, 8'd95};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd108, 8'd105, 8'd87};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd94, 8'd93, 8'd76};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd68};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd63};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd66};
					endcase
				end
				`ybit'd82: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd33};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd32};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd31};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd34};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd33};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd33};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd40};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd40};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd40};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd41};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd49};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd59};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd65};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd52, 8'd59, 8'd72};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd76};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd60, 8'd69, 8'd82};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd85};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd64, 8'd75, 8'd75};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd63, 8'd80, 8'd64};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd68, 8'd84, 8'd57};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd67, 8'd84, 8'd51};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd68, 8'd85, 8'd51};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd48};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd68, 8'd85, 8'd49};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd70, 8'd87, 8'd50};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd70, 8'd87, 8'd51};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd70, 8'd87, 8'd53};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd70, 8'd87, 8'd53};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd69, 8'd86, 8'd52};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd68, 8'd85, 8'd51};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd66, 8'd83, 8'd51};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd67, 8'd80, 8'd49};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd68, 8'd81, 8'd49};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd68, 8'd83, 8'd50};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd70, 8'd83, 8'd51};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd70, 8'd82, 8'd56};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd69, 8'd81, 8'd60};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd69, 8'd80, 8'd64};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd67, 8'd78, 8'd66};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd66, 8'd75, 8'd68};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd60, 8'd69, 8'd80};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd97};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd112};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd122};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd121};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd119};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd115};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd113};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd109};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd109};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd113};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd115};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd114};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd115};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd114};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd115};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd114};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd117};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd48, 8'd54, 8'd112};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd104};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd56, 8'd59, 8'd85};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd61, 8'd62, 8'd62};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd48};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd64, 8'd67, 8'd46};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd64, 8'd63, 8'd45};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd63, 8'd60, 8'd43};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd61, 8'd64, 8'd45};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd47};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd47};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd51};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd53};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd79, 8'd89, 8'd53};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd78, 8'd87, 8'd59};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd76, 8'd83, 8'd74};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd79, 8'd84, 8'd91};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd94, 8'd97, 8'd103};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd115, 8'd112, 8'd105};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd103};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd119, 8'd116, 8'd98};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd93};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd103, 8'd100, 8'd83};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd80};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd84};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd88};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd121, 8'd116, 8'd94};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd123, 8'd117, 8'd96};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd90};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd79};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd94, 8'd91, 8'd76};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd75};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd78};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd87};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd93};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd94};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd93};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd95};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd125, 8'd123, 8'd99};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd131, 8'd128, 8'd103};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd141, 8'd135, 8'd108};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd144, 8'd139, 8'd110};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd111};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd112};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd116};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd144, 8'd138, 8'd114};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd141, 8'd135, 8'd111};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd135, 8'd129, 8'd105};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd126, 8'd124, 8'd101};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd94};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd90};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd80};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd72};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd64};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd64};
					endcase
				end
				`ybit'd83: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd31};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd31};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd31};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd33};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd33};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd34};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd40};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd43};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd49};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd51};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd46, 8'd53, 8'd58};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd57};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd56};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd55};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd58};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd62, 8'd76, 8'd62};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd64, 8'd78, 8'd64};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd65, 8'd80, 8'd66};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd65, 8'd81, 8'd58};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd65, 8'd84, 8'd52};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd68, 8'd85, 8'd48};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd47};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd66, 8'd84, 8'd46};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd48};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd46};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd47};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd69, 8'd87, 8'd48};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd48};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd70, 8'd87, 8'd50};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd68, 8'd87, 8'd49};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd68, 8'd86, 8'd48};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd68, 8'd84, 8'd48};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd67, 8'd83, 8'd47};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd69, 8'd83, 8'd47};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd70, 8'd84, 8'd47};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd71, 8'd85, 8'd48};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd70, 8'd84, 8'd48};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd71, 8'd85, 8'd49};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd70, 8'd83, 8'd52};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd68, 8'd81, 8'd53};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd64, 8'd76, 8'd62};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd79};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd97};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd110};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd120};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd117};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd118};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd112};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd107};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd99};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd98};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd54, 8'd61, 8'd105};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd110};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd113};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd113};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd113};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd113};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd115};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd116};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd115};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd115};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd47, 8'd53, 8'd109};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd95};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd75};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd58, 8'd60, 8'd54};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd59, 8'd64, 8'd44};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd63, 8'd64, 8'd44};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd62, 8'd61, 8'd44};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd61, 8'd57, 8'd41};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd60, 8'd62, 8'd44};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd64, 8'd73, 8'd45};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd45};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd51};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd49};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd49};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd51};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd51};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd76, 8'd88, 8'd53};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd75, 8'd83, 8'd63};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd74, 8'd81, 8'd78};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd84, 8'd87, 8'd93};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd105, 8'd104, 8'd98};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd96};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd91};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd85};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd80};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd78};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd81};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd86};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd120, 8'd115, 8'd94};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd123, 8'd119, 8'd98};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd93};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd84};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd78};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd74};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd75};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd102, 8'd99, 8'd81};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd83};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd82};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd79};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd104, 8'd103, 8'd82};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd93};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd131, 8'd126, 8'd102};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd140, 8'd134, 8'd107};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd109};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd112};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd148, 8'd143, 8'd114};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd146, 8'd140, 8'd115};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd112};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd138, 8'd132, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd134, 8'd128, 8'd104};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd100};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd120, 8'd96};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd93};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd81};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd72};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd64};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd62};
					endcase
				end
				`ybit'd84: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd31};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd31};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd32};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd32};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd31};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd44, 8'd56, 8'd32};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd38};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd45};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd50};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd56};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd62};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd58};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd51};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd50};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd60, 8'd73, 8'd47};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd63, 8'd79, 8'd50};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd66, 8'd82, 8'd53};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd64, 8'd83, 8'd55};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd65, 8'd85, 8'd49};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd67, 8'd84, 8'd48};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd66, 8'd84, 8'd46};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd66, 8'd84, 8'd46};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd68, 8'd82, 8'd46};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd44};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd66, 8'd83, 8'd45};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd67, 8'd81, 8'd45};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd67, 8'd85, 8'd47};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd69, 8'd84, 8'd48};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd70, 8'd84, 8'd48};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd47};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd47};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd71, 8'd84, 8'd48};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd69, 8'd83, 8'd47};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd67, 8'd80, 8'd56};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd60, 8'd72, 8'd67};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd85};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd102};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd110};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd47, 8'd53, 8'd115};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd115};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd46, 8'd53, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd50, 8'd58, 8'd102};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd52, 8'd64, 8'd90};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd85};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd94};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd102};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd104};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd109};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd110};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd108};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd107};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd48, 8'd54, 8'd109};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd47, 8'd53, 8'd109};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd111};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd110};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd109};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd104};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd86};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd65};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd59, 8'd61, 8'd47};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd58, 8'd61, 8'd41};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd63, 8'd62, 8'd44};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd61, 8'd58, 8'd43};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd60, 8'd54, 8'd41};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd58, 8'd59, 8'd42};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd43};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd44};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd47};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd48};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd50};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd47};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd77, 8'd89, 8'd51};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd56};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd73, 8'd80, 8'd69};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd77, 8'd82, 8'd82};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd91, 8'd93, 8'd95};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd94};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd88};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd102, 8'd99, 8'd82};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd76};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd76};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd78};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd102, 8'd99, 8'd80};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd87};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd94};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd93};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd87};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd99, 8'd96, 8'd79};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd73};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd94, 8'd93, 8'd75};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd76};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd76};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd72};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd65};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd68};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd79};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd114, 8'd112, 8'd90};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd131, 8'd125, 8'd102};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd140, 8'd135, 8'd106};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd111};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd113};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd145, 8'd140, 8'd111};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd142, 8'd137, 8'd112};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd140, 8'd134, 8'd110};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd137, 8'd131, 8'd107};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd133, 8'd127, 8'd103};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd126, 8'd123, 8'd98};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd93};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd114, 8'd112, 8'd91};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd81};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd89, 8'd88, 8'd71};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd78, 8'd74, 8'd65};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd62};
					endcase
				end
				`ybit'd85: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd43, 8'd56, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd44, 8'd57, 8'd29};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd44, 8'd57, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd31};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd28};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd29};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd37};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd44};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd52};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd59};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd61};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd51, 8'd63, 8'd55};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd55, 8'd67, 8'd46};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd57, 8'd74, 8'd43};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd61, 8'd78, 8'd45};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd64, 8'd81, 8'd44};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd66, 8'd84, 8'd46};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd45};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd45};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd45};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd45};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd84, 8'd46};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd67, 8'd82, 8'd45};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd66, 8'd80, 8'd44};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd43};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd62, 8'd77, 8'd42};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd43};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd65, 8'd78, 8'd43};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd66, 8'd78, 8'd44};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd66, 8'd80, 8'd45};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd67, 8'd82, 8'd46};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd68, 8'd82, 8'd46};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd70, 8'd84, 8'd47};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd69, 8'd84, 8'd45};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd69, 8'd84, 8'd47};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd68, 8'd83, 8'd43};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd67, 8'd80, 8'd50};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd61, 8'd74, 8'd60};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd76};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd93};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd110};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd118};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd51, 8'd54, 8'd117};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd52, 8'd54, 8'd117};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd119};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd114};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd114};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd98};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd83};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd51, 8'd66, 8'd73};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd85};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd92};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd96};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd102};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd107};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd103};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd101};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd100};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd48, 8'd54, 8'd104};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd104};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd105};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd104};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd99};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd54, 8'd61, 8'd79};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd58, 8'd60, 8'd57};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd59, 8'd58, 8'd43};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd58, 8'd57, 8'd41};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd60, 8'd59, 8'd41};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd60, 8'd56, 8'd44};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd59, 8'd52, 8'd41};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd57, 8'd58, 8'd38};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd42};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd46};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd47};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd49};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd49};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd48};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd52};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd72, 8'd81, 8'd59};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd73, 8'd79, 8'd76};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd90};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd95, 8'd95, 8'd94};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd98, 8'd99, 8'd85};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd96, 8'd94, 8'd79};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd93, 8'd89, 8'd74};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd75};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd76};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd95, 8'd94, 8'd78};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd80};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd107, 8'd106, 8'd86};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd109, 8'd108, 8'd86};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd83};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd76};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd73};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd75};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd75};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd74};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd66};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd59};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd56};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd59};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd69};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd79};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd120, 8'd117, 8'd94};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd134, 8'd128, 8'd105};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd140, 8'd135, 8'd106};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd143, 8'd138, 8'd109};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd142, 8'd136, 8'd112};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd140, 8'd134, 8'd110};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd137, 8'd131, 8'd107};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd134, 8'd128, 8'd104};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd131, 8'd125, 8'd101};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd98};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd95};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd90};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd81};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd70};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd78, 8'd75, 8'd63};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd62};
					endcase
				end
				`ybit'd86: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd43, 8'd56, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd32};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd44, 8'd56, 8'd33};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd32};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd29};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd29};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd35};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd44};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd49};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd52};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd55};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd50};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd59, 8'd72, 8'd45};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd59, 8'd76, 8'd44};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd62, 8'd79, 8'd47};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd63, 8'd80, 8'd44};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd63, 8'd81, 8'd43};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd62, 8'd80, 8'd42};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd64, 8'd82, 8'd44};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd45};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd66, 8'd80, 8'd44};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd65, 8'd78, 8'd46};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd61, 8'd74, 8'd43};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd61, 8'd69, 8'd41};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd60, 8'd68, 8'd42};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd60, 8'd71, 8'd42};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd63, 8'd74, 8'd44};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd64, 8'd78, 8'd43};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd67, 8'd81, 8'd45};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd67, 8'd81, 8'd45};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd68, 8'd82, 8'd46};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd69, 8'd84, 8'd45};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd67, 8'd81, 8'd45};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd66, 8'd80, 8'd44};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd63, 8'd75, 8'd53};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd56, 8'd68, 8'd67};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd89};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd105};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd113};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd52, 8'd53, 8'd117};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd50, 8'd54, 8'd117};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd114};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd114};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd109};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd100};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd85};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd49, 8'd63, 8'd72};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd49, 8'd63, 8'd73};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd79};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd85};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd94};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd100};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd94};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd89};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd87};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd92};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd93};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd95};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd95};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd90};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd68};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd59, 8'd61, 8'd52};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd40};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd56, 8'd54, 8'd39};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd57, 8'd56, 8'd38};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd58, 8'd54, 8'd42};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd59, 8'd51, 8'd40};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd56, 8'd57, 8'd36};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd42};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd66, 8'd77, 8'd42};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd45};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd47};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd47};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd78, 8'd88, 8'd51};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd48};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd49};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd78, 8'd89, 8'd49};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd79, 8'd90, 8'd48};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd51};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd54};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd65};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd76, 8'd82, 8'd81};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd87, 8'd88, 8'd82};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd90, 8'd91, 8'd78};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd72};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd71};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd73};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd74};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd73};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd75};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd80};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd97, 8'd96, 8'd77};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd75};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd87, 8'd84, 8'd69};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd87, 8'd84, 8'd69};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd75};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd77};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd75};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd59};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd54};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd54};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd61};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd72};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd106, 8'd103, 8'd84};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd124, 8'd119, 8'd96};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd100};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd138, 8'd133, 8'd104};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd138, 8'd132, 8'd108};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd135, 8'd129, 8'd105};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd132, 8'd126, 8'd102};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd130, 8'd124, 8'd100};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd128, 8'd122, 8'd98};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd122, 8'd119, 8'd96};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd94};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd90};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd81};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd87, 8'd86, 8'd67};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd64};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd62};
					endcase
				end
				`ybit'd87: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd40, 8'd52, 8'd35};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd40, 8'd51, 8'd34};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd41, 8'd53, 8'd32};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd33};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd36};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd38};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd41};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd47, 8'd61, 8'd48};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd51};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd55, 8'd70, 8'd49};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd57, 8'd73, 8'd44};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd58, 8'd75, 8'd43};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd61, 8'd78, 8'd41};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd61, 8'd79, 8'd41};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd61, 8'd78, 8'd42};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd61, 8'd79, 8'd41};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd62, 8'd79, 8'd42};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd61, 8'd78, 8'd42};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd61, 8'd79, 8'd41};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd61, 8'd78, 8'd42};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd43};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd66, 8'd80, 8'd44};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd66, 8'd80, 8'd44};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd63, 8'd80, 8'd43};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd60, 8'd76, 8'd39};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd58, 8'd67, 8'd39};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd57, 8'd60, 8'd40};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd55, 8'd58, 8'd37};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd56, 8'd62, 8'd40};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd40};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd61, 8'd75, 8'd40};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd64, 8'd78, 8'd42};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd43};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd67, 8'd81, 8'd45};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd44};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd45};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd62, 8'd79, 8'd47};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd58, 8'd71, 8'd58};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd77};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd93};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd108};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd113};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd113};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd116};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd112};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd111};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd102};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd88};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd72};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd63};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd69};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd74};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd81};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd90};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd85};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd51, 8'd63, 8'd79};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd76};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd80};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd83};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd85};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd85};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd78};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd62};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd56, 8'd57, 8'd47};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd56, 8'd53, 8'd38};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd37};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd57, 8'd54, 8'd39};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd59, 8'd50, 8'd39};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd57, 8'd49, 8'd38};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd55, 8'd54, 8'd40};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd60, 8'd65, 8'd39};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd44};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd46};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd77, 8'd87, 8'd50};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd75, 8'd85, 8'd48};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd46};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd46};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd46};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd46};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd47};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd76, 8'd86, 8'd49};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd77, 8'd88, 8'd48};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd77, 8'd88, 8'd48};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd76, 8'd87, 8'd47};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd49};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd57};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd75, 8'd82, 8'd70};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd84, 8'd85, 8'd76};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd77};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd70};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd71};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd72};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd73};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd72};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd72};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd68};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd64};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd60};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd63};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd70};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd77};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd99, 8'd96, 8'd79};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd94, 8'd91, 8'd74};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd68};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd73, 8'd70, 8'd60};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd55};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd57};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd65};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd94, 8'd93, 8'd75};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd108, 8'd107, 8'd83};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd92};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd95};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd122, 8'd121, 8'd94};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd120, 8'd119, 8'd91};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd89};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd120, 8'd114, 8'd89};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd119, 8'd118, 8'd90};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd119, 8'd117, 8'd93};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd93};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd89};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd81};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd69};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd76, 8'd73, 8'd64};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd62};
					endcase
				end
				`ybit'd88: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd41, 8'd52, 8'd33};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd39};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd39};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd41, 8'd52, 8'd37};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd39};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd44};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd45};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd43};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd50, 8'd66, 8'd41};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd54, 8'd70, 8'd45};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd57, 8'd74, 8'd43};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd58, 8'd75, 8'd40};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd60, 8'd78, 8'd40};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd59, 8'd77, 8'd39};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd59, 8'd77, 8'd39};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd59, 8'd76, 8'd40};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd59, 8'd77, 8'd39};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd59, 8'd76, 8'd40};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd59, 8'd77, 8'd40};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd59, 8'd78, 8'd39};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd59, 8'd76, 8'd40};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd41};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd43};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd43};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd61, 8'd77, 8'd41};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd39};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd56, 8'd57, 8'd38};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd54, 8'd50, 8'd39};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd53, 8'd49, 8'd36};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd51, 8'd57, 8'd35};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd60, 8'd74, 8'd39};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd41};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd65, 8'd79, 8'd43};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd41};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd41};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd42};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd59, 8'd74, 8'd47};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd61};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd81};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd44, 8'd51, 8'd96};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd107};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd112};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd113};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd115};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd51, 8'd112};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd100};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd91};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd67};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd65, 8'd57};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd52, 8'd68, 8'd56};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd54, 8'd69, 8'd59};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd65};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd52, 8'd60, 8'd74};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd72};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd66};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd60};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd52, 8'd64, 8'd65};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd68};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd49, 8'd64, 8'd71};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd71};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd64};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd53};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd56, 8'd57, 8'd42};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd37};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd53, 8'd50, 8'd35};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd55, 8'd52, 8'd37};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd56, 8'd48, 8'd37};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd56, 8'd48, 8'd37};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd53, 8'd52, 8'd38};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd58, 8'd63, 8'd37};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd41};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd46};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd46};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd47};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd46};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd44};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd44};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd44};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd73, 8'd84, 8'd44};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd74, 8'd85, 8'd45};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd74, 8'd85, 8'd45};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd73, 8'd83, 8'd49};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd71, 8'd80, 8'd47};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd74, 8'd83, 8'd60};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd84, 8'd87, 8'd66};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd70};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd68};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd65};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd71};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd75};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd75};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd70};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd56};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd52};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd56};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd64};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd75};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd80};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd79};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd95, 8'd94, 8'd76};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd66};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd61};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd58};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd61};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd85, 8'd84, 8'd66};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd74};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd81};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd83};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd82};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd81};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd103, 8'd100, 8'd78};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd106, 8'd99, 8'd79};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd85};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd90};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd91};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd89};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd81};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd67};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd62};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd58};
					endcase
				end
				`ybit'd89: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd50, 8'd36};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd44};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd38};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd36};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd43};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd45};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd41};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd41};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd55, 8'd67, 8'd41};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd55, 8'd71, 8'd42};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd59, 8'd76, 8'd39};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd58, 8'd75, 8'd39};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd58, 8'd75, 8'd39};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd57, 8'd74, 8'd38};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd57, 8'd74, 8'd38};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd56, 8'd73, 8'd37};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd57, 8'd73, 8'd37};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd56, 8'd73, 8'd37};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd58, 8'd74, 8'd38};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd60, 8'd74, 8'd39};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd58, 8'd75, 8'd39};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd61, 8'd75, 8'd39};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd63, 8'd77, 8'd41};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd64, 8'd77, 8'd41};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd60, 8'd76, 8'd39};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd37};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd52, 8'd55, 8'd34};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd48, 8'd35};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd47, 8'd48, 8'd34};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd50, 8'd53, 8'd35};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd37};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd38};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd62, 8'd76, 8'd41};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd62, 8'd76, 8'd40};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd62, 8'd76, 8'd39};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd62, 8'd76, 8'd41};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd60, 8'd74, 8'd41};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd57, 8'd73, 8'd45};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd54, 8'd66, 8'd60};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd78};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd93};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd105};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd91};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd67};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd49};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd47};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd55, 8'd70, 8'd51};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd54};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd59};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd58, 8'd64, 8'd59};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd53};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd50};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd54};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd58};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd52, 8'd68, 8'd57};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd54, 8'd69, 8'd60};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd53, 8'd69, 8'd54};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd45};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd55, 8'd58, 8'd42};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd53, 8'd54, 8'd36};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd51, 8'd52, 8'd34};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd53, 8'd49, 8'd34};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd55, 8'd46, 8'd37};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd52, 8'd43, 8'd36};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd50, 8'd49, 8'd33};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd56, 8'd60, 8'd38};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd64, 8'd73, 8'd44};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd46};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd44};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd44};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd43};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd45};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd43};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd45};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd43};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd46};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd71, 8'd82, 8'd51};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd81, 8'd84, 8'd63};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd85, 8'd86, 8'd68};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd65};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd64};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd66};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd71};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd73};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd74};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd70};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd81, 8'd78, 8'd63};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd56};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd51};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd54};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd60};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd72};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd79};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd87};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd98, 8'd97, 8'd78};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd71};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd62};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd61};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd65};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd67};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd69};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd68};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd66};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd65};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd87, 8'd86, 8'd66};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd74};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd82};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd88};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd88};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd102, 8'd99, 8'd80};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd66};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd60};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
					endcase
				end
				`ybit'd90: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd51, 8'd36};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd43};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd41, 8'd52, 8'd37};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd38};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd40};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd41};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd38};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd40};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd55, 8'd71, 8'd40};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd56, 8'd73, 8'd37};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd56, 8'd73, 8'd38};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd57, 8'd73, 8'd42};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd56, 8'd72, 8'd37};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd55, 8'd72, 8'd37};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd55, 8'd71, 8'd36};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd35};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd56, 8'd72, 8'd37};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd56, 8'd72, 8'd37};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd56, 8'd72, 8'd37};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd59, 8'd74, 8'd38};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd61, 8'd75, 8'd39};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd61, 8'd75, 8'd39};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd58, 8'd73, 8'd38};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd37};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd35};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd50, 8'd49, 8'd34};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd46, 8'd48, 8'd34};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd50, 8'd53, 8'd35};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd37};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd38};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd60, 8'd74, 8'd39};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd61, 8'd75, 8'd39};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd58, 8'd71, 8'd38};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd56, 8'd72, 8'd40};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd55};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd71};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd88};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd110};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd113};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd113};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd113};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd113};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd114};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd111};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd91};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd66};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd47};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd41};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd53, 8'd69, 8'd40};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd41};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd57, 8'd69, 8'd46};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd47};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd62, 8'd70, 8'd42};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd41};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd44};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd52, 8'd68, 8'd44};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd53, 8'd72, 8'd47};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd55, 8'd73, 8'd48};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd52, 8'd71, 8'd41};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd36};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd37};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd54, 8'd56, 8'd37};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd52, 8'd53, 8'd35};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd54, 8'd49, 8'd35};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd53, 8'd45, 8'd35};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd52, 8'd43, 8'd35};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd49, 8'd48, 8'd33};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd53, 8'd57, 8'd35};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd60, 8'd69, 8'd40};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd44};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd44};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd43};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd41};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd42};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd43};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd43};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd46};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd55};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd83, 8'd85, 8'd62};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd64};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd63};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd63};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd73};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd79};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd76};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd70};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd61};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd55};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd55};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd59};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd74};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd109, 8'd106, 8'd85};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd88};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd111, 8'd111, 8'd86};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd79};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd89, 8'd88, 8'd68};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd64};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd63};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd81, 8'd77, 8'd65};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd79, 8'd75, 8'd63};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd75, 8'd72, 8'd60};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd55};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd59};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd67};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd75};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd107, 8'd104, 8'd85};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd87};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd83};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd71};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd64};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
					endcase
				end
				`ybit'd91: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd38, 8'd49, 8'd33};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd39, 8'd50, 8'd36};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd41, 8'd53, 8'd33};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd44, 8'd56, 8'd35};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd38};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd39};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd35};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd37};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd40};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd38};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd40};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd38};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd37};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd40};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd40};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd35};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd34};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd50, 8'd34};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd47, 8'd48, 8'd31};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd51, 8'd53, 8'd35};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd36};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd39};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd36};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd36};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd40};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd58, 8'd71, 8'd41};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd50};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd65};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd85};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd101};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd107};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd48, 8'd49, 8'd113};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd108};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd109};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd110};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd109};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd47, 8'd49, 8'd109};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd108};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd113};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd104};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd42, 8'd49, 8'd91};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd68};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd49, 8'd64, 8'd43};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd37};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd40};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd61, 8'd72, 8'd41};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd59, 8'd72, 8'd41};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd39};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd37};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd52, 8'd68, 8'd38};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd53, 8'd69, 8'd39};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd54, 8'd70, 8'd41};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd51, 8'd67, 8'd38};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd36};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd37};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd37};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd54, 8'd55, 8'd35};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd54, 8'd50, 8'd37};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd53, 8'd46, 8'd33};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd52, 8'd42, 8'd34};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd47, 8'd46, 8'd34};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd35};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd58, 8'd67, 8'd38};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd41};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd41};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd41};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd41};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd44};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd44};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd42};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd44};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd71, 8'd81, 8'd47};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd57};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd81, 8'd84, 8'd62};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd59};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd64};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd92, 8'd91, 8'd71};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd80};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd81};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd75};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd85, 8'd84, 8'd68};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd61};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd58};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd69};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd82};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd92};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd93};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd112, 8'd110, 8'd88};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd79};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd71};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd69};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd64};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd58};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd54};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd49};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd58, 8'd58, 8'd46};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd60, 8'd60, 8'd48};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd66, 8'd63, 8'd52};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd59};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd68};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd78};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd83};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd106, 8'd104, 8'd83};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd100, 8'd99, 8'd79};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd88, 8'd86, 8'd73};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd60};
					endcase
				end
				`ybit'd92: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd28};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd39, 8'd50, 8'd31};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd32};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd34};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd35};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd36};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd34};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd35};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd34};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd36};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd36};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd53, 8'd67, 8'd33};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd54, 8'd67, 8'd37};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd38};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd38};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd37};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd34};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd52, 8'd64, 8'd34};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd35};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd35};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd53, 8'd67, 8'd35};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd32};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd33};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd47, 8'd48, 8'd33};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd46, 8'd33};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd49, 8'd51, 8'd35};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd35};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd36};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd36};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd36};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd37};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd59, 8'd72, 8'd37};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd58, 8'd71, 8'd43};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd51};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd69};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd85};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd101};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd106};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd109};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd109};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd112};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd109};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd108};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd108};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd109};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd109};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd108};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd108};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd104};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd46, 8'd49, 8'd106};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd106};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd111};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd109};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd102};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd90};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd67};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd43};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd35};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd50, 8'd65, 8'd36};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd37};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd59, 8'd72, 8'd37};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd57, 8'd74, 8'd38};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd53, 8'd69, 8'd36};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd50, 8'd67, 8'd35};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd50, 8'd67, 8'd34};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd50, 8'd67, 8'd35};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd51, 8'd66, 8'd35};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd37};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd33};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd34};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd37};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd35};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd54, 8'd50, 8'd36};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd54, 8'd45, 8'd33};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd50, 8'd40, 8'd32};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd45, 8'd44, 8'd32};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd49, 8'd52, 8'd33};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd37};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd39};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd39};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd40};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd39};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd41};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd42};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd69, 8'd78, 8'd43};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd75, 8'd81, 8'd49};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd81, 8'd84, 8'd61};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd65};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd63};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd61};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd69};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd77};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd82};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd101, 8'd98, 8'd79};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd91, 8'd90, 8'd71};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd64};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd59};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd58};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd62};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd85, 8'd82, 8'd66};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd77};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd93};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd121, 8'd117, 8'd93};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd116, 8'd112, 8'd88};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd83};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd77};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd72};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd62};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd71, 8'd68, 8'd57};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd63, 8'd60, 8'd51};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd45};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd45};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd62, 8'd59, 8'd52};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd55};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd62};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd87, 8'd85, 8'd72};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd99, 8'd96, 8'd77};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd82};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd82};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd77};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd88, 8'd85, 8'd68};
					endcase
				end
				`ybit'd93: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd27};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd40, 8'd51, 8'd27};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd43, 8'd56, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd32};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd34};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd34};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd34};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd33};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd35};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd35};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd38};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd34};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd33};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd33};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd34};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd34};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd33};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd32};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd48, 8'd32};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd45, 8'd43, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd46, 8'd44, 8'd31};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd32};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd33};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd36};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd59, 8'd73, 8'd40};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd57, 8'd69, 8'd45};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd61};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd45, 8'd52, 8'd77};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd40, 8'd46, 8'd93};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd102};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd107};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd109};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd102};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd102};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd103};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd107};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd111};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd109};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd103};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd91};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd69};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd43};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd48, 8'd64, 8'd35};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd49, 8'd63, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd55, 8'd69, 8'd34};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd54, 8'd71, 8'd35};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd50, 8'd67, 8'd35};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd49, 8'd66, 8'd34};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd49, 8'd66, 8'd34};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd49, 8'd66, 8'd34};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd50, 8'd65, 8'd32};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd34};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd33};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd33};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd35};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd35};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd53, 8'd50, 8'd35};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd51, 8'd43, 8'd31};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd49, 8'd40, 8'd31};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd44, 8'd43, 8'd31};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd48, 8'd50, 8'd32};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd35};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd41};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd39};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd43};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd71, 8'd78, 8'd45};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd80, 8'd85, 8'd56};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd86, 8'd86, 8'd65};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd66};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd66};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd71};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd76};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd74};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd89, 8'd87, 8'd69};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd64};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd57};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd59};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd82, 8'd79, 8'd64};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd71};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd79};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd113, 8'd111, 8'd88};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd124, 8'd118, 8'd94};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd125, 8'd119, 8'd95};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd90};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd111, 8'd109, 8'd86};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd101, 8'd100, 8'd79};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd90, 8'd89, 8'd69};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd63};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd55};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd48};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd46};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd60, 8'd57, 8'd50};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd50};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd79, 8'd76, 8'd63};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd70};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd76};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd105, 8'd103, 8'd82};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd103, 8'd101, 8'd80};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd74};
					endcase
				end
				`ybit'd94: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd25};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd28};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd32};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd33};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd35};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd33};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd34};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd34};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd34};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd34};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd37};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd33};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd33};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd31};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd32};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd50, 8'd52, 8'd31};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd50, 8'd48, 8'd28};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd50, 8'd53, 8'd32};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd32};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd32};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd29};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd46, 8'd43, 8'd32};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd42, 8'd39, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd43, 8'd41, 8'd29};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd45, 8'd47, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd33};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd36};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd37};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd58, 8'd71, 8'd41};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd56, 8'd70, 8'd40};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd52, 8'd66, 8'd50};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd70};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd40, 8'd48, 8'd86};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd99};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd106};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd106};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd43, 8'd46, 8'd109};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd43, 8'd46, 8'd109};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd105};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd105};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd105};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd105};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd105};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd106};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd106};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd106};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd107};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd43, 8'd46, 8'd110};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd104};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd100};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd99};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd100};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd106};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd43, 8'd46, 8'd108};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd110};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd106};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd106};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd103};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd88};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd63};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd44};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd50, 8'd67, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd48, 8'd65, 8'd33};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd48, 8'd62, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd34};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd52, 8'd64, 8'd35};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd51, 8'd68, 8'd36};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd51, 8'd68, 8'd36};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd48, 8'd64, 8'd32};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd48, 8'd64, 8'd35};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd35};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd35};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd32};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd31};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd33};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd33};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd33};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd50, 8'd48, 8'd33};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd46, 8'd44, 8'd31};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd49, 8'd39, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd44, 8'd41, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd45, 8'd47, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd52, 8'd56, 8'd34};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd58, 8'd67, 8'd38};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd39};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd38};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd38};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd40};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd39};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd42};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd69, 8'd79, 8'd42};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd38};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd40};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd67, 8'd78, 8'd42};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd74, 8'd84, 8'd50};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd86, 8'd88, 8'd64};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd84, 8'd85, 8'd68};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd80, 8'd77, 8'd63};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd61};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd85, 8'd82, 8'd63};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd89, 8'd85, 8'd67};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd85, 8'd84, 8'd64};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd61};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd55};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd67, 8'd66, 8'd50};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd58};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd78, 8'd75, 8'd60};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd66};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd91, 8'd90, 8'd72};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd81};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd115, 8'd113, 8'd90};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd124, 8'd122, 8'd99};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd127, 8'd121, 8'd97};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd120, 8'd118, 8'd95};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd113, 8'd110, 8'd87};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd104, 8'd101, 8'd79};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd75};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd65};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd72, 8'd69, 8'd59};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd63, 8'd60, 8'd50};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd47};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd59, 8'd59, 8'd47};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd52};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd63};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd69};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd105, 8'd102, 8'd83};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd78};
					endcase
				end
				`ybit'd95: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd27};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd29};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd33};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd35};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd37};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd52, 8'd66, 8'd31};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd36};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd36};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd35};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd34};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd34};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd35};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd32};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd47, 8'd49, 8'd32};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd48, 8'd44, 8'd31};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd51, 8'd43, 8'd32};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd49, 8'd48, 8'd34};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd33};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd31};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd27};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd45, 8'd41, 8'd29};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd29};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd46, 8'd49, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd31};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd33};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd33};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd34};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd57, 8'd71, 8'd36};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd55, 8'd69, 8'd39};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd46};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd61};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd82};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd37, 8'd43, 8'd95};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd102};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd107};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd109};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd109};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd109};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd104};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd42, 8'd45, 8'd109};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd42, 8'd45, 8'd109};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd109};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd105};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd100};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd44, 8'd51, 8'd96};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd90};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd44, 8'd51, 8'd91};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd98};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd41, 8'd47, 8'd103};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd105};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd99};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd44, 8'd51, 8'd84};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd51, 8'd59, 8'd59};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd42};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd51, 8'd69, 8'd32};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd51, 8'd68, 8'd36};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd48, 8'd62, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd32};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd33};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd49, 8'd66, 8'd34};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd48, 8'd65, 8'd33};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd47, 8'd64, 8'd32};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd46, 8'd62, 8'd33};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd33};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd32};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd31};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd32};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd32};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd32};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd49, 8'd46, 8'd31};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd46, 8'd43, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd47, 8'd37, 8'd28};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd44, 8'd40, 8'd29};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd43, 8'd45, 8'd28};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd32};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd35};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd40};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd38};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd60, 8'd69, 8'd39};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd39};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd42};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd72, 8'd82, 8'd48};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd82, 8'd84, 8'd60};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd83, 8'd84, 8'd67};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd77, 8'd79, 8'd68};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd78, 8'd75, 8'd64};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd79, 8'd75, 8'd62};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd78, 8'd75, 8'd62};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd58};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd67, 8'd64, 8'd54};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd64, 8'd61, 8'd50};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd48};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd56};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd77, 8'd74, 8'd59};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd81, 8'd78, 8'd63};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd86, 8'd85, 8'd66};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd73};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd107, 8'd105, 8'd81};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd93};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd125, 8'd119, 8'd95};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd96};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd116, 8'd114, 8'd91};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd110, 8'd108, 8'd85};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd101, 8'd99, 8'd79};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd71};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd67};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd55};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd50};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd60, 8'd60, 8'd48};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd48};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd56};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd66};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd71};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd81};
					endcase
				end
				`ybit'd96: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd26};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd28};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd32};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd35};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd35};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd36};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd53, 8'd67, 8'd32};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd53, 8'd67, 8'd31};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd52, 8'd66, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd35};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd35};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd34};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd33};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd32};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd44, 8'd47, 8'd28};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd27};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd44, 8'd40, 8'd29};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd46, 8'd40, 8'd28};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd45, 8'd45, 8'd31};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd29};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd31};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd50, 8'd34};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd46, 8'd48, 8'd33};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd45, 8'd46, 8'd31};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd32};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd33};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd34};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd33};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd33};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd42};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd61, 8'd50};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd70};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd38, 8'd45, 8'd90};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd98};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd104};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd104};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd44, 8'd46, 8'd104};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd100};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd90};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd86};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd82};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd80};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd90};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd97};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd45, 8'd47, 8'd103};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd46, 8'd100};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd44, 8'd46, 8'd100};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd93};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd77};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd53};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd40};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd51, 8'd68, 8'd33};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd49, 8'd66, 8'd34};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd32};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd32};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd33};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd46, 8'd63, 8'd31};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd46, 8'd63, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd46, 8'd63, 8'd31};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd45, 8'd61, 8'd32};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd46, 8'd61, 8'd32};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd33};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd31};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd29};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd31};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd46, 8'd44, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd43, 8'd41, 8'd29};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd45, 8'd36, 8'd31};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd45, 8'd36, 8'd31};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd27};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd33};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd36};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd35};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd35};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd64, 8'd76, 8'd40};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd38};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd41};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd64, 8'd76, 8'd40};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd40};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd68, 8'd78, 8'd41};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd40};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd67, 8'd77, 8'd43};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd75, 8'd80, 8'd52};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd77, 8'd79, 8'd65};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd74, 8'd75, 8'd70};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd73, 8'd73, 8'd67};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd77, 8'd73, 8'd64};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd76, 8'd73, 8'd58};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd46};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd54, 8'd53, 8'd45};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd54, 8'd54, 8'd46};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd62, 8'd59, 8'd52};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd61};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd80, 8'd77, 8'd64};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd64};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd69};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd73};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd109, 8'd107, 8'd83};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd114, 8'd112, 8'd88};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd117, 8'd111, 8'd88};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd112, 8'd109, 8'd86};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd108, 8'd106, 8'd82};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd104, 8'd102, 8'd81};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd74};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd68};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd61, 8'd61, 8'd49};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd62, 8'd62, 8'd50};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd58};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd64};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd71};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
					endcase
				end
				`ybit'd97: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd29};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd31};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd32};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd31};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd32};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd32};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd32};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd33};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd33};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd33};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd53, 8'd68, 8'd33};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd35};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd33};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd31};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd46, 8'd43, 8'd31};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd44, 8'd40, 8'd28};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd44, 8'd36, 8'd28};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd41, 8'd38, 8'd27};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd44, 8'd39, 8'd27};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd44, 8'd45, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd31};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd29};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd32};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd33};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd54, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd33};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd33};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd51, 8'd59, 8'd35};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd32};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd33};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd35};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd35};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd47};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd62};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd38, 8'd46, 8'd81};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd35, 8'd40, 8'd95};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd35, 8'd39, 8'd101};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd36, 8'd40, 8'd103};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd106};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd106};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd106};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd108};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd40, 8'd43, 8'd106};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd107};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd102};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd104};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd102};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd40, 8'd46, 8'd103};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd44, 8'd46, 8'd98};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd86};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd76};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd51, 8'd57, 8'd72};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd50, 8'd57, 8'd65};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd66};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd75};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd82};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd85};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd88};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd88};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd45, 8'd52, 8'd82};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd67};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd46};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd34};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd49, 8'd66, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd46, 8'd63, 8'd31};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd31};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd45, 8'd62, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd46, 8'd63, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd46, 8'd62, 8'd31};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd45, 8'd61, 8'd32};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd43, 8'd58, 8'd29};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd31};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd29};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd29};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd29};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd29};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd28};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd43, 8'd40, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd44, 8'd35, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd44, 8'd35, 8'd29};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd26};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd31};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd36};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd35};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd62, 8'd74, 8'd38};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd37};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd61, 8'd73, 8'd37};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd37};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd37};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd36};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd39};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd39};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd64, 8'd75, 8'd45};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd66, 8'd74, 8'd58};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd65, 8'd69, 8'd73};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd68, 8'd71, 8'd75};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd77, 8'd74, 8'd70};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd63};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd45};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd51, 8'd51, 8'd43};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd51, 8'd52, 8'd43};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd58, 8'd55, 8'd48};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd58};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd62};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd62};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd85, 8'd82, 8'd65};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd68};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd75};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd101, 8'd97, 8'd79};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd104, 8'd97, 8'd79};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd99, 8'd95, 8'd76};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd96, 8'd93, 8'd74};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd96, 8'd94, 8'd73};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd99, 8'd98, 8'd76};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd73};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd81, 8'd80, 8'd60};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd63, 8'd62, 8'd50};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd61, 8'd62, 8'd49};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd51};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd77, 8'd74, 8'd57};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd63};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd70};
					endcase
				end
				`ybit'd98: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd33};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd33};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd31};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd29};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd29};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd31};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd32};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd32};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd51, 8'd64, 8'd34};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd52, 8'd64, 8'd34};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd34};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd34};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd31};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd33};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd46, 8'd49, 8'd28};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd46, 8'd44, 8'd28};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd44, 8'd41, 8'd28};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd42, 8'd38, 8'd26};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd40, 8'd36, 8'd25};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd40, 8'd36, 8'd25};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd40, 8'd41, 8'd28};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd43, 8'd46, 8'd25};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd31};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd33};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd32};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd32};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd33};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd29};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd32};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd29};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd31};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd50, 8'd55, 8'd32};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd39};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd51};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd40, 8'd48, 8'd67};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd35, 8'd41, 8'd84};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd33, 8'd38, 8'd95};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd35, 8'd40, 8'd97};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd36, 8'd41, 8'd98};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd38, 8'd42, 8'd103};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd105};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd105};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd101};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd107};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd107};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd103};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd103};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd107};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd107};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd106};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd41, 8'd44, 8'd98};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd91};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd51, 8'd54, 8'd74};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd54, 8'd59, 8'd61};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd56};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd55};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd52};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd57};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd63};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd65};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd70};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd46, 8'd53, 8'd68};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd47, 8'd53, 8'd66};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd54};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd41};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd32};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd45, 8'd62, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd44, 8'd59, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd42, 8'd58, 8'd29};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd44, 8'd60, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd44, 8'd60, 8'd31};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd44, 8'd57, 8'd29};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd32};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd45, 8'd52, 8'd28};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd27};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd28};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd28};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd27};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd31};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd40, 8'd41, 8'd29};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd41, 8'd36, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd43, 8'd34, 8'd29};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd43, 8'd34, 8'd29};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd41, 8'd39, 8'd27};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd46, 8'd48, 8'd29};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd36};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd36};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd36};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd36};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd36};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd38};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd35};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd40};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd59, 8'd65, 8'd56};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd58, 8'd62, 8'd69};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd61, 8'd65, 8'd76};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd74, 8'd73, 8'd74};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd81, 8'd78, 8'd67};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd61};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd51};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd54, 8'd54, 8'd46};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd51, 8'd51, 8'd43};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd56, 8'd53, 8'd46};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd49};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd59};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd63};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd64};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd85, 8'd82, 8'd65};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd66};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd65};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd64};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd62};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd65};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd72};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd77};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd76};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd70};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd61};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd48};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd52};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd58};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd64};
					endcase
				end
				`ybit'd99: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd33};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd32};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd28};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd27};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd28};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd29};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd47, 8'd61, 8'd31};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd33};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd51, 8'd63, 8'd33};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd33};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd32};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd28};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd46, 8'd43, 8'd27};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd45, 8'd40, 8'd29};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd45, 8'd38, 8'd27};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd43, 8'd37, 8'd25};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd42, 8'd37, 8'd28};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd40, 8'd41, 8'd29};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd40, 8'd46, 8'd29};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd28};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd29};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd33};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd32};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd31};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd29};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd32};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd28};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd31};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd47, 8'd48, 8'd29};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd31};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd33};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd38};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd57};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd39, 8'd46, 8'd74};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd35, 8'd42, 8'd84};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd35, 8'd40, 8'd93};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd36, 8'd41, 8'd94};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd95};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd98};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd99};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd100};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd101};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd102};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd102};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd102};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd103};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd103};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd103};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd105};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd105};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd102};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd102};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd39, 8'd42, 8'd103};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd104};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd105};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd104};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd41, 8'd44, 8'd95};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd83};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd62};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd47};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd58, 8'd65, 8'd41};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd39};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd38};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd42};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd44};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd53, 8'd60, 8'd47};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd51};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd51, 8'd57, 8'd51};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd48};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd42};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd35};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd27};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd29};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd44, 8'd61, 8'd29};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd29};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd29};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd28};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd27};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd27};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd27};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd27};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd39, 8'd40, 8'd27};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd41, 8'd36, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd43, 8'd35, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd42, 8'd34, 8'd29};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd39, 8'd37, 8'd25};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd45, 8'd47, 8'd28};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd34};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd60, 8'd69, 8'd34};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd36};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd35};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd35};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd39};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd38};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd38};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd36};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd36};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd34};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd56, 8'd63, 8'd48};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd54, 8'd58, 8'd64};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd75};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd70, 8'd69, 8'd77};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd82, 8'd78, 8'd72};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd67};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd60};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd61, 8'd60, 8'd50};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd45};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd56, 8'd53, 8'd45};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd47};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd51};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd57};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd63};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd64};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd62};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd60};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd58};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd52};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd51};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd56};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd82, 8'd78, 8'd66};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd72};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd98, 8'd97, 8'd75};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd72};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd67};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd62};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd70, 8'd67, 8'd54};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd50};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd57};
					endcase
				end
				`ybit'd100: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd52, 8'd66, 8'd32};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd52, 8'd66, 8'd31};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd49, 8'd63, 8'd28};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd27};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd28};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd29};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd29};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd27};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd42, 8'd42, 8'd28};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd43, 8'd39, 8'd27};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd43, 8'd39, 8'd28};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd43, 8'd39, 8'd27};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd44, 8'd39, 8'd26};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd28};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd44, 8'd46, 8'd29};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd27};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd29};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd32};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd34};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd29};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd29};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd44, 8'd46, 8'd29};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd44, 8'd45, 8'd29};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd45, 8'd48, 8'd31};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd34};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd49};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd62};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd40, 8'd47, 8'd71};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd40, 8'd46, 8'd77};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd80};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd41, 8'd47, 8'd81};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd85};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd40, 8'd46, 8'd85};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd42, 8'd45, 8'd92};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd42, 8'd45, 8'd93};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd39, 8'd45, 8'd94};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd38, 8'd44, 8'd94};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd39, 8'd45, 8'd96};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd97};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd96};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd97};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd99};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd39, 8'd42, 8'd99};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd98};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd36, 8'd42, 8'd99};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd101};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd100};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd100};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd100};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd39, 8'd46, 8'd92};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd77};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd54, 8'd60, 8'd54};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd39};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd57, 8'd65, 8'd35};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd34};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd34};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd34};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd36};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd55, 8'd63, 8'd37};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd38};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd39};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd38};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd34};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd33};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd27};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd29};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd44, 8'd61, 8'd29};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd42, 8'd59, 8'd29};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd42, 8'd58, 8'd29};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd44, 8'd57, 8'd29};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd28};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd26};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd38, 8'd44, 8'd24};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd37, 8'd38, 8'd25};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd38, 8'd34, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd42, 8'd33, 8'd28};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd43, 8'd34, 8'd28};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd39, 8'd36, 8'd25};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd41, 8'd43, 8'd27};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd51, 8'd57, 8'd31};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd59, 8'd66, 8'd33};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd35};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd35};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd65, 8'd75, 8'd38};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd35};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd36};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd58, 8'd66, 8'd42};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd53, 8'd60, 8'd55};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd55, 8'd60, 8'd68};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd63, 8'd66, 8'd78};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd78};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd88, 8'd85, 8'd74};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd67};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd72, 8'd71, 8'd54};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd47};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd43};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd45};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd56};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd80, 8'd77, 8'd62};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd63};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd63};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd60};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd47};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd43};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd56, 8'd54, 8'd42};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd47};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd55};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd65};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd95, 8'd93, 8'd71};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd76};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd73};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd66};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd76, 8'd73, 8'd56};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd51};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd52};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
					endcase
				end
				`ybit'd101: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd54, 8'd68, 8'd32};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd52, 8'd65, 8'd28};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd28};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd26};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd41, 8'd44, 8'd24};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd41, 8'd42, 8'd28};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd43, 8'd44, 8'd29};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd27};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd28};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd29};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd26};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd26};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd43, 8'd42, 8'd28};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd41, 8'd39, 8'd27};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd44, 8'd38, 8'd27};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd43, 8'd39, 8'd27};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd28};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd44, 8'd43, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd44, 8'd47, 8'd29};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd46, 8'd53, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd34};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd29};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd49, 8'd63, 8'd29};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd26};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd29};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd45, 8'd46, 8'd29};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd46, 8'd46, 8'd29};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd45, 8'd49, 8'd29};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd48, 8'd53, 8'd33};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd44};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd50};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd57};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd58};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd62};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd66};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd45, 8'd52, 8'd66};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd70};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd43, 8'd50, 8'd76};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd79};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd80};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd84};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd87};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd43, 8'd45, 8'd86};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd89};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd41, 8'd45, 8'd90};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd40, 8'd43, 8'd95};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd40, 8'd43, 8'd98};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd94};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd41, 8'd97};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd39, 8'd42, 8'd96};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd39, 8'd41, 8'd98};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd39, 8'd41, 8'd98};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd38, 8'd41, 8'd98};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd41, 8'd46, 8'd87};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd68};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd47};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd37};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd32};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd31};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd44, 8'd59, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd47, 8'd61, 8'd32};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd32};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd31};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd45, 8'd59, 8'd29};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd46, 8'd60, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd46, 8'd60, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd42, 8'd50, 8'd27};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd41, 8'd48, 8'd28};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd25};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd22};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd36, 8'd37, 8'd25};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd36, 8'd34, 8'd23};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd41, 8'd32, 8'd24};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd41, 8'd32, 8'd24};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd38, 8'd35, 8'd23};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd40, 8'd39, 8'd24};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd28};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd31};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd33};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd33};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd35};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd33};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd35};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd35};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd35};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd57, 8'd64, 8'd32};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd57, 8'd65, 8'd32};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd35};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd36};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd36};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd61, 8'd70, 8'd41};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd57, 8'd66, 8'd48};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd55, 8'd61, 8'd60};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd58, 8'd61, 8'd78};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd70, 8'd74, 8'd81};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd89, 8'd85, 8'd77};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd74};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd66};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd70, 8'd67, 8'd55};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd61, 8'd58, 8'd49};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd44};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd48};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd60};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd63};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd66};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd63};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd58};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd64, 8'd61, 8'd52};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd43};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd41};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd43};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd48};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd60};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd87, 8'd86, 8'd66};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd98, 8'd95, 8'd75};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd76};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd71};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd63};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd73, 8'd72, 8'd55};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd50};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
					endcase
				end
				`ybit'd102: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd52, 8'd66, 8'd31};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd27};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd27};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd41, 8'd44, 8'd26};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd42, 8'd38, 8'd26};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd38, 8'd26};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd44, 8'd39, 8'd27};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd44, 8'd42, 8'd27};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd28};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd27};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd40, 8'd48, 8'd25};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd39, 8'd42, 8'd26};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd40, 8'd37, 8'd25};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd41, 8'd39, 8'd26};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd43, 8'd42, 8'd25};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd43, 8'd45, 8'd27};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd26};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd46, 8'd50, 8'd29};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd33};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd29};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd29};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd49, 8'd63, 8'd28};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd29};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd46, 8'd53, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd29};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd49, 8'd54, 8'd29};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd32};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd37};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd36};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd41};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd42};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd43};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd46};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd47};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd52};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd54};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd58};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd58};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd49, 8'd53, 8'd63};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd65};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd45, 8'd50, 8'd67};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd43, 8'd50, 8'd71};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd72};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd43, 8'd50, 8'd78};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd81};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd40, 8'd47, 8'd78};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd83};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd86};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd88};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd87};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd40, 8'd44, 8'd88};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd41, 8'd48, 8'd76};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd47, 8'd53, 8'd60};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd52, 8'd59, 8'd42};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd31};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd31};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd29};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd31};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd50, 8'd64, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd50, 8'd63, 8'd33};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd48, 8'd62, 8'd28};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd28};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd28};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd25};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd40, 8'd48, 8'd25};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd25};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd38, 8'd44, 8'd24};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd35, 8'd36, 8'd23};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd37, 8'd35, 8'd23};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd41, 8'd32, 8'd23};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd41, 8'd32, 8'd23};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd36, 8'd33, 8'd21};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd38, 8'd37, 8'd22};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd26};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd52, 8'd59, 8'd29};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd33};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd35};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd35};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd35};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd31};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd31};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd64, 8'd74, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd66, 8'd77, 8'd35};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd37};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd60, 8'd71, 8'd42};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd52};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd56, 8'd61, 8'd70};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd64, 8'd68, 8'd81};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd81, 8'd81, 8'd81};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd78};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd69};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd59};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd51};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd46};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd45};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd50};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd80, 8'd77, 8'd60};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd88, 8'd85, 8'd68};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd69};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd62};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd58};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd50};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd44};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd56, 8'd54, 8'd42};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd44};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd59};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd69};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd98, 8'd96, 8'd75};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd99, 8'd97, 8'd76};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd68};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd81, 8'd80, 8'd62};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd54};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd51};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
					endcase
				end
				`ybit'd103: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd28};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd41, 8'd54, 8'd24};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd23};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd39, 8'd38, 8'd23};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd39, 8'd35, 8'd24};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd34, 8'd25};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd44, 8'd35, 8'd26};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd43, 8'd39, 8'd27};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd42, 8'd44, 8'd28};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd40, 8'd43, 8'd27};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd37, 8'd39, 8'd24};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd38, 8'd38, 8'd28};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd41, 8'd42, 8'd26};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd45, 8'd47, 8'd28};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd27};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd48, 8'd54, 8'd29};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd31};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd51, 8'd65, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd49, 8'd62, 8'd28};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd45, 8'd59, 8'd29};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd31};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd33};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd33};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd34};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd35};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd35};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd37};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd37};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd40};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd42};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd51, 8'd59, 8'd46};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd47};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd48};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd50};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd54};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd55};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd58};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd60};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd64};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd42, 8'd50, 8'd67};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd42, 8'd49, 8'd71};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd71};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd72};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd73};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd65};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd51, 8'd55, 8'd52};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd51, 8'd59, 8'd37};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd27};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd27};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd54, 8'd66, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd58, 8'd70, 8'd34};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd56, 8'd68, 8'd32};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd50, 8'd65, 8'd34};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd33};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd33};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd54, 8'd66, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd51, 8'd59, 8'd31};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd31};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd29};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd28};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd28};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd24};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd25};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd37, 8'd38, 8'd24};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd37, 8'd35, 8'd25};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd37, 8'd35, 8'd25};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd40, 8'd34, 8'd25};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd36, 8'd39, 8'd22};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd27};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd51, 8'd56, 8'd29};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd33};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd35};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd34};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd33};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd33};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd34};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd62, 8'd72, 8'd35};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd37};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd63, 8'd73, 8'd36};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd37};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd57, 8'd66, 8'd47};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd62};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd57, 8'd62, 8'd80};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd75, 8'd75, 8'd81};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd91, 8'd89, 8'd81};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd97, 8'd93, 8'd74};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd68};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd77, 8'd73, 8'd62};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd50};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd59, 8'd58, 8'd45};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd46};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd51};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd75, 8'd73, 8'd60};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd85, 8'd82, 8'd63};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd69};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd92, 8'd89, 8'd70};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd67};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd60};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd51};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd45};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd44};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd63};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd71};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd74};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd70};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd66};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd57};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd52};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
					endcase
				end
				`ybit'd104: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd27};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd38, 8'd45, 8'd22};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd38, 8'd37, 8'd23};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd39, 8'd31, 8'd23};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd40, 8'd30, 8'd21};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd41, 8'd32, 8'd23};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd41, 8'd33, 8'd23};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd39, 8'd36, 8'd23};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd40, 8'd42, 8'd26};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd40, 8'd48, 8'd25};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd40, 8'd47, 8'd25};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd28};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd40, 8'd43, 8'd22};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd26};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd26};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd27};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd26};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd46, 8'd59, 8'd27};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd47, 8'd61, 8'd28};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd62, 8'd27};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd48, 8'd62, 8'd27};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd31};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd47, 8'd60, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd53, 8'd61, 8'd32};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd33};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd29};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd32};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd33};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd33};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd33};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd48, 8'd61, 8'd35};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd36};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd37};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd39};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd40};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd43};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd47};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd47, 8'd52, 8'd51};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd53};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd54};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd55};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd48};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd40};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd32};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd25};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd28};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd28};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd56, 8'd68, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd59, 8'd72, 8'd36};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd57, 8'd70, 8'd34};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd59, 8'd71, 8'd33};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd57, 8'd69, 8'd33};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd28};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd27};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd24};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd42, 8'd44, 8'd24};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd25};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd26};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd41, 8'd41, 8'd25};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd41, 8'd43, 8'd27};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd28};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd29};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd32};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd33};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd34};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd34};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd37};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd51};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd53, 8'd61, 8'd68};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd63, 8'd68, 8'd80};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd82, 8'd83, 8'd85};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd97, 8'd93, 8'd82};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd69};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd88, 8'd84, 8'd66};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd56};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd62, 8'd61, 8'd49};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd46};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd47};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd53};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd58};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd90, 8'd87, 8'd68};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd95, 8'd92, 8'd73};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd71};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd85, 8'd84, 8'd65};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd73, 8'd73, 8'd54};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd51};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd48};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd55};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd77, 8'd77, 8'd58};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd87, 8'd84, 8'd68};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd67};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd65};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd81, 8'd78, 8'd61};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd54};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd47};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
					endcase
				end
				`ybit'd105: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd38, 8'd45, 8'd22};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd37, 8'd36, 8'd18};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd34, 8'd33, 8'd21};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd35, 8'd30, 8'd19};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd38, 8'd29, 8'd24};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd38, 8'd29, 8'd20};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd39, 8'd31, 8'd22};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd39, 8'd36, 8'd22};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd38, 8'd42, 8'd27};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd38, 8'd48, 8'd24};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd26};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd41, 8'd48, 8'd27};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd39, 8'd46, 8'd25};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd26};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd29};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd29};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd28};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd28};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd45, 8'd58, 8'd28};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd32};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd27};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd32};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd31};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd35};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd34};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd35};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd47, 8'd54, 8'd38};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd38};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd42};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd42};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd40};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd51, 8'd59, 8'd34};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd29};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd55, 8'd67, 8'd31};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd56, 8'd69, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd34};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd56, 8'd65, 8'd32};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd32};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd29};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd26};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd29};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd29};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd47, 8'd50, 8'd28};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd46, 8'd49, 8'd27};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd25};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd26};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd56, 8'd64, 8'd35};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd54, 8'd62, 8'd43};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd62};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd57, 8'd60, 8'd78};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd72, 8'd73, 8'd79};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd91, 8'd90, 8'd80};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd102, 8'd98, 8'd77};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd75};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd65};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd47};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd48};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd51};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd55};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd65};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd93, 8'd91, 8'd70};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd97, 8'd95, 8'd74};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd91, 8'd88, 8'd69};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd61};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd72, 8'd71, 8'd53};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd50};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd48};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd75, 8'd72, 8'd57};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd58};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd60};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd77, 8'd76, 8'd57};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd51};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd50};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd45};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd46};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd46};
					endcase
				end
				`ybit'd106: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd35, 8'd36, 8'd21};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd34, 8'd32, 8'd20};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd33, 8'd31, 8'd23};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd36, 8'd30, 8'd20};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd36, 8'd28, 8'd22};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd34, 8'd30, 8'd20};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd35, 8'd33, 8'd22};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd35, 8'd38, 8'd22};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd39, 8'd43, 8'd22};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd25};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd39, 8'd50, 8'd25};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd38, 8'd52, 8'd24};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd39, 8'd53, 8'd25};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd43, 8'd55, 8'd25};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd41, 8'd59, 8'd27};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd42, 8'd58, 8'd29};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd43, 8'd56, 8'd26};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd44, 8'd57, 8'd27};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd44, 8'd57, 8'd27};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd26};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd27};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd29};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd27};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd27};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd28};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd28};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd25};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd26};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd26};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd27};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd27};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd28};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd27};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd50, 8'd58, 8'd29};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd33};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd28};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd29};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd27};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd56, 8'd68, 8'd32};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd34};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd32};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd29};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd32};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd29};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd25};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd28};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd50, 8'd58, 8'd28};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd28};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd29};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd33};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd31};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd31};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd31};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd28};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd33};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd32};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd32};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd35};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd52, 8'd58, 8'd50};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd53, 8'd56, 8'd70};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd60, 8'd64, 8'd78};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd82, 8'd81, 8'd82};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd99, 8'd94, 8'd82};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd100, 8'd97, 8'd78};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd89, 8'd88, 8'd67};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd61};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd50};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd47};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd47};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd68, 8'd67, 8'd50};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd78, 8'd76, 8'd58};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd87, 8'd84, 8'd64};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd69};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd90, 8'd88, 8'd68};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd62};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd74, 8'd73, 8'd56};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd51};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd49};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd75, 8'd72, 8'd57};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd58};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd44};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd53, 8'd52, 8'd39};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd40};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd56, 8'd54, 8'd41};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd43};
					endcase
				end
				`ybit'd107: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd32, 8'd33, 8'd19};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd35, 8'd33, 8'd21};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd35, 8'd33, 8'd21};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd35, 8'd32, 8'd20};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd36, 8'd32, 8'd22};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd34, 8'd31, 8'd21};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd35, 8'd33, 8'd23};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd34, 8'd41, 8'd22};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd22};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd37, 8'd52, 8'd23};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd38, 8'd52, 8'd24};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd38, 8'd54, 8'd25};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd40, 8'd54, 8'd23};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd41, 8'd57, 8'd26};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd40, 8'd57, 8'd25};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd40, 8'd57, 8'd25};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd39, 8'd56, 8'd25};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd41, 8'd54, 8'd25};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd43, 8'd55, 8'd25};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd29};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd31};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd43, 8'd56, 8'd26};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd42, 8'd55, 8'd25};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd27};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd42, 8'd55, 8'd25};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd26};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd27};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd25};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd41, 8'd47, 8'd23};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd42, 8'd43, 8'd23};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd43, 8'd45, 8'd24};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd25};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd26};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd27};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd28};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd32};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd33};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd34};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd53, 8'd62, 8'd31};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd51, 8'd57, 8'd29};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd53, 8'd61, 8'd27};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd55, 8'd62, 8'd29};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd32};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd33};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd33};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd28};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd28};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd55, 8'd64, 8'd32};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd53, 8'd59, 8'd42};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd59};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd52, 8'd57, 8'd71};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd70, 8'd70, 8'd83};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd89, 8'd86, 8'd83};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd97, 8'd94, 8'd79};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd93, 8'd92, 8'd76};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd66};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd54};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd48};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd46};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd49};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd55};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd76, 8'd59};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd62};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd62};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd76, 8'd75, 8'd58};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd55};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd48};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd50};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd56};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd52};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd47};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd39};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd48, 8'd46, 8'd34};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd44, 8'd44, 8'd32};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd47, 8'd45, 8'd37};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd52, 8'd49, 8'd41};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd56, 8'd54, 8'd42};
					endcase
				end
				`ybit'd108: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd36, 8'd36, 8'd23};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd38, 8'd39, 8'd21};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd39, 8'd40, 8'd21};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd38, 8'd39, 8'd21};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd37, 8'd38, 8'd22};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd33, 8'd36, 8'd20};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd36, 8'd40, 8'd24};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd35, 8'd44, 8'd23};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd35, 8'd50, 8'd22};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd35, 8'd52, 8'd23};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd37, 8'd53, 8'd23};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd39, 8'd55, 8'd25};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd39, 8'd55, 8'd25};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd37, 8'd54, 8'd24};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd37, 8'd53, 8'd24};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd39, 8'd54, 8'd25};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd40, 8'd55, 8'd26};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd42, 8'd55, 8'd25};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd25};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd23};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd27};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd28};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd27};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd24};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd41, 8'd54, 8'd24};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd26};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd43, 8'd55, 8'd25};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd26};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd25};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd23};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd40, 8'd38, 8'd23};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd42, 8'd39, 8'd24};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd42, 8'd47, 8'd24};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd26};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd24};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd27};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd28};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd26};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd26};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd26};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd31};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd32};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd60, 8'd70, 8'd32};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd32};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd29};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd31};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd32};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd49, 8'd56, 8'd28};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd29};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd29};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd29};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd29};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd27};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd27};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd26};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd25};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd29};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd61, 8'd71, 8'd32};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd32};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd29};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd28};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd28};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd53, 8'd61, 8'd34};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd50, 8'd57, 8'd49};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd66};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd60, 8'd60, 8'd81};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd83};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd83, 8'd82, 8'd82};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd84, 8'd83, 8'd76};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd70};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd68, 8'd67, 8'd60};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd63, 8'd62, 8'd50};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd61, 8'd61, 8'd48};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd65, 8'd64, 8'd49};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd52};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd71, 8'd67, 8'd54};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd53};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd50};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd63, 8'd62, 8'd46};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd59, 8'd59, 8'd46};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd44};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd46};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd52};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd54};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd52};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd45};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd51, 8'd49, 8'd36};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd44, 8'd43, 8'd31};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd40, 8'd40, 8'd32};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd42, 8'd41, 8'd34};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd47, 8'd46, 8'd38};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd40};
					endcase
				end
				`ybit'd109: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd38, 8'd42, 8'd24};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd42, 8'd49, 8'd24};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd24};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd43, 8'd51, 8'd25};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd40, 8'd47, 8'd24};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd23};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd24};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd23};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd38, 8'd54, 8'd25};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd42, 8'd55, 8'd25};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd28};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd27};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd27};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd41, 8'd53, 8'd23};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd40, 8'd53, 8'd23};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd24};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd39, 8'd38, 8'd21};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd36, 8'd34, 8'd20};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd39, 8'd37, 8'd22};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd25};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd25};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd28};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd62, 8'd73, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd61, 8'd72, 8'd32};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd28};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd29};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd53, 8'd65, 8'd27};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd49, 8'd55, 8'd27};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd50, 8'd56, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd26};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd31};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd25};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd28};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd31};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd27};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd27};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd33};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd39};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd55};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd50, 8'd53, 8'd74};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd57, 8'd60, 8'd84};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd64, 8'd66, 8'd84};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd66, 8'd67, 8'd80};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd63, 8'd65, 8'd75};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd59, 8'd61, 8'd72};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd59, 8'd59, 8'd61};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd63, 8'd62, 8'd56};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd67, 8'd66, 8'd51};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd70, 8'd68, 8'd53};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd66, 8'd63, 8'd48};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd46};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd40};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd50, 8'd48, 8'd36};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd48, 8'd48, 8'd36};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd53, 8'd51, 8'd38};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd42};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd66, 8'd64, 8'd49};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd73, 8'd72, 8'd54};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd55};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd39};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd45, 8'd45, 8'd33};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd40, 8'd40, 8'd32};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd40, 8'd40, 8'd32};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd44, 8'd44, 8'd35};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd51, 8'd49, 8'd37};
					endcase
				end
				`ybit'd110: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd26};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd23};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd26};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd26};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd24};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd40, 8'd53, 8'd23};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd37, 8'd53, 8'd24};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd33, 8'd52, 8'd22};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd32, 8'd48, 8'd19};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd37, 8'd50, 8'd22};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd39, 8'd53, 8'd24};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd24};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd26};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd23};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd41, 8'd53, 8'd23};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd40, 8'd53, 8'd25};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd25};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd42, 8'd56, 8'd27};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd23};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd40, 8'd41, 8'd22};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd38, 8'd34, 8'd22};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd37, 8'd31, 8'd21};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd39, 8'd18};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd24};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd25};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd27};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd27};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd26};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd32};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd62, 8'd73, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd60, 8'd71, 8'd31};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd29};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd26};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd28};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd26};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd28};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd27};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd29};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd27};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd27};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd27};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd35};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd47, 8'd53, 8'd47};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd64};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd84};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd85};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd83};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd47, 8'd51, 8'd83};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd76};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd51, 8'd53, 8'd68};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd62, 8'd62, 8'd66};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd57};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd52};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd51};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd45};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd50, 8'd50, 8'd37};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd43, 8'd44, 8'd32};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd43, 8'd43, 8'd35};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd45, 8'd45, 8'd33};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd53, 8'd51, 8'd39};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd47};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd71, 8'd69, 8'd53};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd77, 8'd76, 8'd57};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd54};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd47};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd53, 8'd50, 8'd42};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd45, 8'd43, 8'd31};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd42, 8'd39, 8'd31};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd45, 8'd42, 8'd35};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd48, 8'd45, 8'd38};
					endcase
				end
				`ybit'd111: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd26};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd26};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd44, 8'd61, 8'd24};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd44, 8'd60, 8'd24};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd41, 8'd58, 8'd22};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd42, 8'd58, 8'd23};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd42, 8'd55, 8'd25};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd38, 8'd54, 8'd25};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd32, 8'd51, 8'd21};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd19};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd35, 8'd51, 8'd22};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd39, 8'd52, 8'd24};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd42, 8'd55, 8'd27};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd27};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd26};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd49, 8'd57, 8'd29};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd29};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd28};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd27};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd40, 8'd53, 8'd25};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd23};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd23};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd39, 8'd52, 8'd24};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd41, 8'd48, 8'd21};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd36, 8'd38, 8'd18};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd35, 8'd31, 8'd19};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd37, 8'd31, 8'd21};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd37, 8'd39, 8'd18};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd43, 8'd48, 8'd22};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd22};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd23};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd41, 8'd51, 8'd24};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd27};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd27};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd54, 8'd63, 8'd28};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd26};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd25};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd59, 8'd69, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd58, 8'd68, 8'd31};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd28};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd26};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd26};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd29};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd47, 8'd55, 8'd38};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd40, 8'd51, 8'd56};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd38, 8'd45, 8'd75};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd35, 8'd42, 8'd85};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd33, 8'd39, 8'd86};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd34, 8'd40, 8'd89};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd35, 8'd42, 8'd84};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd42, 8'd46, 8'd79};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd55, 8'd58, 8'd71};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd63};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd61};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd74, 8'd72, 8'd57};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd49};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd53, 8'd52, 8'd40};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd44, 8'd44, 8'd33};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd40, 8'd40, 8'd32};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd44, 8'd44, 8'd31};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd51, 8'd49, 8'd36};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd43};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd68, 8'd66, 8'd49};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd75, 8'd74, 8'd56};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd60};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd72, 8'd71, 8'd55};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd48};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd40};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd47, 8'd45, 8'd37};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd45, 8'd42, 8'd35};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd47, 8'd44, 8'd37};
					endcase
				end
				`ybit'd112: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd22};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd46, 8'd60, 8'd25};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd46, 8'd60, 8'd25};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd46, 8'd60, 8'd25};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd43, 8'd60, 8'd24};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd41, 8'd58, 8'd22};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd39, 8'd56, 8'd21};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd38, 8'd55, 8'd23};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd36, 8'd53, 8'd21};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd31, 8'd48, 8'd18};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd31, 8'd50, 8'd20};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd31, 8'd50, 8'd20};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd35, 8'd50, 8'd21};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd39, 8'd52, 8'd23};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd21};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd41, 8'd49, 8'd25};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd36, 8'd47, 8'd19};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd36, 8'd47, 8'd19};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd36, 8'd44, 8'd20};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd38, 8'd46, 8'd22};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd38, 8'd48, 8'd21};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd23};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd23};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd38, 8'd49, 8'd20};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd38, 8'd41, 8'd21};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd36, 8'd33, 8'd17};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd34, 8'd32, 8'd19};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd35, 8'd35, 8'd21};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd35, 8'd42, 8'd19};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd42, 8'd48, 8'd22};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd23};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd24};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd38, 8'd48, 8'd21};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd38, 8'd48, 8'd21};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd25};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd26};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd25};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd25};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd24};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd24};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd26};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd28};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd29};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd29};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd51, 8'd63, 8'd27};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd29};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd27};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd24};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd48, 8'd56, 8'd33};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd47};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd64};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd32, 8'd39, 8'd81};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd28, 8'd35, 8'd86};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd28, 8'd35, 8'd88};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd29, 8'd35, 8'd87};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd33, 8'd41, 8'd81};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd49, 8'd51, 8'd77};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd65, 8'd65, 8'd67};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd63};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd60};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd56};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd46};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd51, 8'd48, 8'd40};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd42, 8'd42, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd46, 8'd43, 8'd36};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd50, 8'd47, 8'd36};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd41};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd48};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd72, 8'd71, 8'd53};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd58};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd58};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd56};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd63, 8'd60, 8'd49};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd53, 8'd51, 8'd39};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd47, 8'd45, 8'd33};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd46, 8'd44, 8'd32};
					endcase
				end
				`ybit'd113: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd44, 8'd58, 8'd23};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd44, 8'd58, 8'd23};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd43, 8'd57, 8'd22};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd40, 8'd57, 8'd21};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd38, 8'd55, 8'd19};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd36, 8'd53, 8'd18};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd34, 8'd51, 8'd19};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd33, 8'd50, 8'd18};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd32, 8'd48, 8'd19};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd32, 8'd48, 8'd19};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd30, 8'd49, 8'd19};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd31, 8'd50, 8'd20};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd34, 8'd50, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd23};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd25};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd43, 8'd57, 8'd22};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd50, 8'd61, 8'd27};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd26};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd26};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd39, 8'd47, 8'd23};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd36, 8'd42, 8'd20};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd35, 8'd41, 8'd18};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd19};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd35, 8'd44, 8'd20};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd34, 8'd44, 8'd20};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd33, 8'd35, 8'd20};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd33, 8'd29, 8'd18};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd32, 8'd31, 8'd18};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd35, 8'd35, 8'd21};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd37, 8'd43, 8'd21};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd23};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd44, 8'd52, 8'd24};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd40, 8'd51, 8'd20};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd38, 8'd48, 8'd21};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd24};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd25};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd27};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd25};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd22};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd23};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd25};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd44, 8'd50, 8'd24};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd24};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd25};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd26};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd27};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd28};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd29};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd29};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd25};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd27};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd50, 8'd59, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd26};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd29};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd46, 8'd54, 8'd38};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd38, 8'd49, 8'd54};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd33, 8'd41, 8'd74};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd28, 8'd36, 8'd86};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd27, 8'd33, 8'd90};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd27, 8'd33, 8'd91};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd29, 8'd35, 8'd87};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd82};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd55, 8'd59, 8'd70};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd74, 8'd74, 8'd69};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd63};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd79, 8'd78, 8'd58};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd70, 8'd69, 8'd49};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd43};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd48, 8'd48, 8'd36};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd48, 8'd44, 8'd38};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd48, 8'd46, 8'd34};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd52, 8'd50, 8'd38};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd44};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd68, 8'd67, 8'd49};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd76, 8'd75, 8'd55};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd59};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd57};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd73, 8'd71, 8'd55};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd63, 8'd61, 8'd48};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd52, 8'd50, 8'd38};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd47, 8'd45, 8'd34};
					endcase
				end
				`ybit'd114: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd42, 8'd56, 8'd21};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd41, 8'd55, 8'd20};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd41, 8'd55, 8'd20};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd41, 8'd55, 8'd20};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd38, 8'd55, 8'd19};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd36, 8'd53, 8'd21};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd34, 8'd51, 8'd19};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd33, 8'd50, 8'd18};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd32, 8'd48, 8'd19};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd31, 8'd47, 8'd18};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd38, 8'd51, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd40, 8'd53, 8'd22};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd26};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd22};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd19};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd35, 8'd36, 8'd19};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd34, 8'd35, 8'd18};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd34, 8'd38, 8'd19};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd35, 8'd40, 8'd18};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd20};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd19};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd36, 8'd44, 8'd20};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd34, 8'd42, 8'd19};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd32, 8'd38, 8'd16};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd32, 8'd31, 8'd18};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd15};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd33, 8'd29, 8'd17};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd33, 8'd37, 8'd20};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd42, 8'd19};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd20};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd24};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd24};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd40, 8'd50, 8'd23};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd23};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd27};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd21};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd22};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd28};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd51, 8'd60, 8'd26};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd55, 8'd67, 8'd29};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd29};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd27};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd22};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd28};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd51, 8'd58, 8'd33};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd44};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd65};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd31, 8'd38, 8'd80};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd27, 8'd34, 8'd88};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd26, 8'd32, 8'd87};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd27, 8'd34, 8'd89};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd34, 8'd38, 8'd82};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd48, 8'd49, 8'd78};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd71};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd79, 8'd79, 8'd68};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd82, 8'd80, 8'd65};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd57};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd52};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd42};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd50, 8'd48, 8'd36};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd49, 8'd47, 8'd35};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd51, 8'd49, 8'd38};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd53, 8'd54, 8'd40};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd62, 8'd60, 8'd45};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd70, 8'd69, 8'd51};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd77, 8'd76, 8'd58};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd82, 8'd79, 8'd60};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd61};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd55};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd44};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd51, 8'd49, 8'd36};
					endcase
				end
				`ybit'd115: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd53, 8'd19};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd39, 8'd52, 8'd20};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd37, 8'd51, 8'd19};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd37, 8'd51, 8'd19};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd36, 8'd52, 8'd20};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd34, 8'd51, 8'd19};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd32, 8'd49, 8'd17};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd31, 8'd47, 8'd16};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd31, 8'd47, 8'd18};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd31, 8'd47, 8'd18};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd38, 8'd51, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd41, 8'd54, 8'd23};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd22};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd25};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd25};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd23};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd25};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd21};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd39, 8'd47, 8'd19};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd37, 8'd36, 8'd18};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd34, 8'd30, 8'd18};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd34, 8'd30, 8'd19};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd35, 8'd34, 8'd20};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd35, 8'd40, 8'd18};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd19};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd34, 8'd42, 8'd18};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd19};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd32, 8'd40, 8'd16};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd30, 8'd34, 8'd13};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd30, 8'd28, 8'd15};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd29, 8'd27, 8'd14};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd33, 8'd30, 8'd17};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd33, 8'd37, 8'd19};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd44, 8'd18};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd25};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd41, 8'd52, 8'd22};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd39, 8'd50, 8'd21};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd20};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd22};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd25};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd47, 8'd56, 8'd26};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd23};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd21};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd26};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd26};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd48, 8'd57, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd22};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd22};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd27};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd56, 8'd67, 8'd28};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd27};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd23};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd24};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd23};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd25};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd51, 8'd62, 8'd27};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd27};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd56, 8'd66, 8'd29};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd59, 8'd70, 8'd29};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd58, 8'd69, 8'd28};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd27};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd27};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd27};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd24};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd24};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd21};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd21};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd24};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd28};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd38};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd43, 8'd49, 8'd56};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd35, 8'd42, 8'd72};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd28, 8'd34, 8'd86};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd26, 8'd32, 8'd89};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd27, 8'd33, 8'd88};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd28, 8'd35, 8'd87};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd38, 8'd42, 8'd81};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd55, 8'd55, 8'd75};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd73, 8'd72, 8'd69};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd66};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd81, 8'd80, 8'd60};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd72, 8'd70, 8'd56};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd63, 8'd60, 8'd47};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd41};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd50, 8'd48, 8'd37};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd51, 8'd48, 8'd37};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd51, 8'd52, 8'd38};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd41};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd65, 8'd63, 8'd47};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd73, 8'd72, 8'd53};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd81, 8'd79, 8'd61};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd64};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd80, 8'd78, 8'd59};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd48};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd58, 8'd56, 8'd44};
					endcase
				end
				`ybit'd116: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd38, 8'd51, 8'd21};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd36, 8'd49, 8'd21};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd34, 8'd47, 8'd19};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd34, 8'd47, 8'd19};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd36, 8'd49, 8'd19};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd33, 8'd50, 8'd17};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd31, 8'd48, 8'd17};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd19};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd20};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd40, 8'd52, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd24};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd48, 8'd59, 8'd24};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd23};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd22};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd24};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd48, 8'd60, 8'd24};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd23};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd37, 8'd41, 8'd19};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd33, 8'd31, 8'd17};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd31, 8'd27, 8'd16};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd31, 8'd27, 8'd16};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd33, 8'd32, 8'd18};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd34, 8'd38, 8'd17};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd18};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd36, 8'd44, 8'd20};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd34, 8'd42, 8'd18};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd32, 8'd40, 8'd17};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd32, 8'd35, 8'd14};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd33, 8'd29, 8'd17};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd31, 8'd29, 8'd16};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd34, 8'd32, 8'd18};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd34, 8'd38, 8'd19};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd44, 8'd19};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd41, 8'd52, 8'd22};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd39, 8'd50, 8'd20};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd35, 8'd45, 8'd18};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd37, 8'd48, 8'd21};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd23};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd26};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd45, 8'd53, 8'd24};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd23};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd55, 8'd65, 8'd28};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd23};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd22};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd26};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd57, 8'd68, 8'd28};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd55, 8'd66, 8'd26};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd54, 8'd64, 8'd27};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd23};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd22};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd50, 8'd62, 8'd26};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd32};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd48, 8'd55, 8'd48};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd40, 8'd47, 8'd64};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd30, 8'd40, 8'd79};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd27, 8'd34, 8'd87};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd26, 8'd33, 8'd88};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd27, 8'd32, 8'd88};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd31, 8'd38, 8'd85};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd79};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd60, 8'd63, 8'd72};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd75, 8'd74, 8'd70};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd77, 8'd76, 8'd68};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd71, 8'd70, 8'd63};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd63, 8'd62, 8'd57};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd55, 8'd54, 8'd50};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd50, 8'd49, 8'd44};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd48, 8'd47, 8'd41};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd49, 8'd49, 8'd37};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd40};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd60, 8'd58, 8'd45};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd67, 8'd66, 8'd47};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd78, 8'd77, 8'd59};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd86, 8'd83, 8'd64};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd84, 8'd81, 8'd62};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd79, 8'd77, 8'd57};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd69, 8'd67, 8'd52};
					endcase
				end
				`ybit'd117: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd37, 8'd50, 8'd20};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd35, 8'd48, 8'd20};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd32, 8'd45, 8'd17};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd33, 8'd46, 8'd18};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd34, 8'd47, 8'd19};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd18};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd32, 8'd48, 8'd16};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd28, 8'd44, 8'd16};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd31, 8'd47, 8'd18};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd34, 8'd47, 8'd20};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd40, 8'd52, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd24};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd22};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd22};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd22};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd22};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd22};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd22};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd22};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd23};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd24};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd23};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd47, 8'd59, 8'd23};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd19};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd19};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd32, 8'd34, 8'd14};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd30, 8'd27, 8'd16};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd30, 8'd22, 8'd16};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd32, 8'd24, 8'd18};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd32, 8'd30, 8'd17};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd34, 8'd37, 8'd20};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd34, 8'd42, 8'd18};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd36, 8'd44, 8'd20};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd36, 8'd44, 8'd20};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd19};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd35, 8'd39, 8'd19};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd33, 8'd37, 8'd19};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd33, 8'd36, 8'd19};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd32, 8'd36, 8'd19};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd35, 8'd41, 8'd18};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd39, 8'd44, 8'd21};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd19};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd38, 8'd48, 8'd21};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd24};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd22};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd21};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd24};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd26};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd26};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd21};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd24};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd49, 8'd58, 8'd24};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd24};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd23};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd54, 8'd65, 8'd24};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd22};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd22};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd22};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd24};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd23};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd23};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd23};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd25};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd53, 8'd64, 8'd28};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd38};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd53};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd33, 8'd43, 8'd71};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd29, 8'd36, 8'd86};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd26, 8'd32, 8'd88};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd27, 8'd32, 8'd88};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd28, 8'd35, 8'd87};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd34, 8'd40, 8'd83};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd48, 8'd52, 8'd78};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd60, 8'd61, 8'd74};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd65, 8'd64, 8'd72};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd62, 8'd61, 8'd68};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd55, 8'd56, 8'd62};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd50, 8'd51, 8'd59};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd46, 8'd47, 8'd52};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd45, 8'd47, 8'd42};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd46, 8'd48, 8'd36};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd50, 8'd50, 8'd38};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd57, 8'd55, 8'd42};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd48};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd72, 8'd71, 8'd54};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd81, 8'd80, 8'd60};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd63};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd85, 8'd83, 8'd61};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd76, 8'd74, 8'd56};
					endcase
				end
				`ybit'd118: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd37, 8'd50, 8'd20};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd36, 8'd49, 8'd20};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd32, 8'd45, 8'd17};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd32, 8'd45, 8'd17};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd33, 8'd46, 8'd18};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd33, 8'd50, 8'd18};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd32, 8'd49, 8'd17};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd36, 8'd49, 8'd21};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd40, 8'd51, 8'd22};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd25};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd20};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd45, 8'd56, 8'd22};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd22};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd22};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd23};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd23};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd46, 8'd58, 8'd22};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd45, 8'd57, 8'd21};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd19};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd32, 8'd40, 8'd17};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd28, 8'd30, 8'd15};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd27, 8'd24, 8'd13};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd30, 8'd21, 8'd16};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd32, 8'd23, 8'd18};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd32, 8'd30, 8'd16};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd33, 8'd35, 8'd18};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd34, 8'd43, 8'd19};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd36, 8'd44, 8'd20};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd37, 8'd45, 8'd21};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd37, 8'd45, 8'd21};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd20};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd37, 8'd42, 8'd20};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd39, 8'd42, 8'd20};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd20};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd38, 8'd43, 8'd20};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd40, 8'd45, 8'd22};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd36, 8'd46, 8'd19};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd39, 8'd49, 8'd22};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd24};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd51, 8'd61, 8'd26};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd25};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd24};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd22};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd46, 8'd57, 8'd22};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd42, 8'd52, 8'd18};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd23};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd22};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd21};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd21};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd22};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd21};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd22};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd22};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd53, 8'd63, 8'd27};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd52, 8'd62, 8'd31};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd50, 8'd57, 8'd45};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd38, 8'd50, 8'd64};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd33, 8'd41, 8'd79};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd29, 8'd35, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd28, 8'd33, 8'd89};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd27, 8'd32, 8'd89};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd31, 8'd37, 8'd87};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd36, 8'd43, 8'd81};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd44, 8'd48, 8'd79};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd44, 8'd49, 8'd78};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd43, 8'd47, 8'd76};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd41, 8'd44, 8'd74};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd39, 8'd42, 8'd68};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd37, 8'd40, 8'd61};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd38, 8'd42, 8'd51};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd44, 8'd44, 8'd42};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd48, 8'd47, 8'd41};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd54, 8'd52, 8'd39};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd59, 8'd57, 8'd44};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd66, 8'd65, 8'd48};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd75, 8'd74, 8'd54};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd60};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd86, 8'd84, 8'd62};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd81, 8'd78, 8'd60};
					endcase
				end
				`ybit'd119: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd39, 8'd52, 8'd22};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd37, 8'd50, 8'd19};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd32, 8'd45, 8'd15};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd32, 8'd45, 8'd17};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd34, 8'd47, 8'd19};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd33, 8'd49, 8'd18};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd33, 8'd50, 8'd18};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd34, 8'd51, 8'd19};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd35, 8'd48, 8'd18};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd31, 8'd47, 8'd18};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd30, 8'd46, 8'd17};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd35, 8'd48, 8'd18};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd42, 8'd54, 8'd19};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd42, 8'd53, 8'd19};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd19};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd19};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd44, 8'd55, 8'd21};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd19};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd18};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd30, 8'd33, 8'd13};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd27, 8'd25, 8'd14};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd25, 8'd20, 8'd15};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd25, 8'd21, 8'd14};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd27, 8'd22, 8'd16};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd26, 8'd28, 8'd13};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd31, 8'd35, 8'd18};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd32, 8'd41, 8'd17};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd35, 8'd43, 8'd19};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd36, 8'd45, 8'd18};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd36, 8'd45, 8'd18};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd37, 8'd47, 8'd20};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd19};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd19};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd18};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd18};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd36, 8'd45, 8'd18};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd19};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd25};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd19};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd20};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd44, 8'd53, 8'd24};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd45, 8'd54, 8'd25};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd21};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd21};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd45, 8'd51, 8'd23};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd46, 8'd52, 8'd23};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd46, 8'd56, 8'd22};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd49, 8'd59, 8'd24};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd25};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd48, 8'd58, 8'd23};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd20};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd43, 8'd52, 8'd23};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd18};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd21};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd23};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd47, 8'd57, 8'd22};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd42, 8'd51, 8'd22};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd43, 8'd53, 8'd20};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd45, 8'd55, 8'd21};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd44, 8'd54, 8'd20};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd21};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd21};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd41, 8'd50, 8'd21};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd19};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd39, 8'd48, 8'd19};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd19};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd37, 8'd46, 8'd19};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd38, 8'd47, 8'd20};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd40, 8'd49, 8'd20};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd46, 8'd55, 8'd21};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd49, 8'd60, 8'd24};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd52, 8'd61, 8'd39};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd43, 8'd54, 8'd52};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd37, 8'd44, 8'd74};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd31, 8'd38, 8'd86};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd28, 8'd34, 8'd87};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd28, 8'd35, 8'd89};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd28, 8'd35, 8'd89};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd28, 8'd36, 8'd83};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd28, 8'd37, 8'd82};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd30, 8'd37, 8'd82};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd27, 8'd34, 8'd80};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd27, 8'd34, 8'd80};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd27, 8'd34, 8'd77};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd29, 8'd35, 8'd73};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd35, 8'd37, 8'd63};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd37, 8'd40, 8'd48};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd44, 8'd44, 8'd39};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd51, 8'd50, 8'd37};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd55, 8'd53, 8'd41};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd61, 8'd59, 8'd46};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd67, 8'd65, 8'd50};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd76, 8'd73, 8'd54};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd83, 8'd80, 8'd61};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd84, 8'd82, 8'd61};
					endcase
				end
			endcase
		end
	end

endmodule