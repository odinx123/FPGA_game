module showMap(clk, rst, X, Y, mapR, mapG, mapB);

	parameter xbit = 10, ybit = 9;
	input clk, rst;
	input [xbit-1:0] X;
	input [ybit-1:0] Y;
	output [7:0] mapR, mapG, mapB;
	reg [7:0] mapR, mapG, mapB;

	always @(posedge clk) begin
		if(!rst) begin
			mapR <= 8'd255;
			mapG <= 8'd255;
			mapB <= 8'd255;
		end
		else begin
			case(Y)
				`ybit'd0: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd1: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd217};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd2: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd3: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd4: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd89};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd91};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd218, 8'd217, 8'd215};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd91};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd218, 8'd216, 8'd219};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd89};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd5: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd254, 8'd254, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd216};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd216};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd253, 8'd254, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd216};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd216};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd216, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd6: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd7: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd8: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd184, 8'd124, 8'd81};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd252};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd85};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd253};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd219, 8'd215, 8'd220};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd85};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd219, 8'd217, 8'd214};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd184, 8'd124, 8'd81};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd9: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd216, 8'd216};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd254};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd254};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd88};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd180, 8'd124, 8'd88};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd249};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd183, 8'd122, 8'd90};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd250};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd10: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd251};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd90};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd87};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd181, 8'd124, 8'd87};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd88};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd11: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd218, 8'd217, 8'd215};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd121, 8'd92};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd90};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd12: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd121, 8'd92};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd90};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd216, 8'd219};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd215};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd183, 8'd125, 8'd79};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd13: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd216};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd84};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd251};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd83};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd91};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd250};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd14: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd251};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd187, 8'd122, 8'd83};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd86};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd86};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd86};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd250};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd15: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd16: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd17: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd215, 8'd217, 8'd219};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd253};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd253};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd90};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd18: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd121, 8'd90};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd85};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd19: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd213};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd20: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd251};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd21: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd213};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd22: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd23: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd24: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd25: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd26: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd89};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd90};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd218, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd215};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd214};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd85};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd218, 8'd216, 8'd218};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd218, 8'd216, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd90};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd218, 8'd216, 8'd219};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd89};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd27: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd215};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd184, 8'd122, 8'd91};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd28: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd90};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd29: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd90};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd182, 8'd123, 8'd89};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd88};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd181, 8'd124, 8'd87};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd30: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd250};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd179, 8'd124, 8'd89};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd253};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd89};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd251};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd218, 8'd217, 8'd215};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd218, 8'd217, 8'd215};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd215, 8'd219, 8'd212};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd31: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd214, 8'd218, 8'd221};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd32: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd214, 8'd218, 8'd221};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd33: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd214, 8'd218, 8'd221};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd252};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd91};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd183, 8'd122, 8'd91};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd87};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd187, 8'd121, 8'd87};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd34: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd88};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd86};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd90};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd35: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd121, 8'd92};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd90};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd36: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd121, 8'd92};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd218};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd183, 8'd122, 8'd92};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd37: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd220, 8'd215, 8'd215};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd121, 8'd92};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd219};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd88};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd253};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd184, 8'd124, 8'd84};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd86};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd38: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd90};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd253};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd88};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd186, 8'd122, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd39: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd85};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd214, 8'd218, 8'd219};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd215};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd253, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd85};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd40: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd41: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd42: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd218, 8'd216};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd43: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd89};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd216};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd254};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd89};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd254};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd44: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd215};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd220, 8'd216, 8'd215};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd219};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd253};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd218, 8'd216, 8'd217};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd253};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd45: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd46: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd255};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd217};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd255};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd216, 8'd217, 8'd218};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
				`ybit'd47: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd185, 8'd123, 8'd86};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd87};
					endcase
				end
			endcase
		end
	end

endmodule