module wall(clk, rst, X, Y, is_wall);

	parameter xbit = 10, ybit = 9;
	input clk, rst;
	input [xbit-1:0] X;
	input [ybit-1:0] Y;
	output reg is_wall;

	always @(posedge clk, negedge rst) begin
		if(!rst) begin
		is_wall <= 1'b0;
		end
		else begin
			case(Y)
				`ybit'd0: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b0;
						`xbit'd2: is_wall <= 1'b0;
						`xbit'd3: is_wall <= 1'b0;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b0;
						`xbit'd6: is_wall <= 1'b0;
						`xbit'd7: is_wall <= 1'b0;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b0;
						`xbit'd10: is_wall <= 1'b0;
						`xbit'd11: is_wall <= 1'b0;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b0;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b0;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b0;
						`xbit'd26: is_wall <= 1'b0;
						`xbit'd27: is_wall <= 1'b0;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b0;
						`xbit'd30: is_wall <= 1'b0;
						`xbit'd31: is_wall <= 1'b0;
						`xbit'd32: is_wall <= 1'b0;
						`xbit'd33: is_wall <= 1'b0;
						`xbit'd34: is_wall <= 1'b0;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b0;
						`xbit'd37: is_wall <= 1'b0;
						`xbit'd38: is_wall <= 1'b0;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b0;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b0;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b0;
						`xbit'd53: is_wall <= 1'b0;
						`xbit'd54: is_wall <= 1'b0;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b0;
						`xbit'd57: is_wall <= 1'b0;
						`xbit'd58: is_wall <= 1'b0;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b0;
						`xbit'd61: is_wall <= 1'b0;
						`xbit'd62: is_wall <= 1'b0;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd1: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd2: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd3: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd4: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b0;
						`xbit'd10: is_wall <= 1'b0;
						`xbit'd11: is_wall <= 1'b0;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b0;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b0;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b0;
						`xbit'd26: is_wall <= 1'b0;
						`xbit'd27: is_wall <= 1'b0;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b0;
						`xbit'd37: is_wall <= 1'b0;
						`xbit'd38: is_wall <= 1'b0;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b0;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b0;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b0;
						`xbit'd53: is_wall <= 1'b0;
						`xbit'd54: is_wall <= 1'b0;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd5: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd6: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd7: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd8: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd9: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd10: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd11: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd12: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd13: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd14: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd15: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd16: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd17: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd18: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b0;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd19: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd20: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd21: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b0;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b0;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b0;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd22: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd23: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd24: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd25: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd26: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b0;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b0;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b0;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd27: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd28: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd29: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b0;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd30: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd31: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd32: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd33: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd34: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd35: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd36: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd37: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd38: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd39: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd40: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd41: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd42: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd43: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b0;
						`xbit'd10: is_wall <= 1'b0;
						`xbit'd11: is_wall <= 1'b0;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b0;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b0;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b0;
						`xbit'd26: is_wall <= 1'b0;
						`xbit'd27: is_wall <= 1'b0;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b0;
						`xbit'd37: is_wall <= 1'b0;
						`xbit'd38: is_wall <= 1'b0;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b0;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b0;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b0;
						`xbit'd53: is_wall <= 1'b0;
						`xbit'd54: is_wall <= 1'b0;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd44: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd45: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd46: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b1;
						`xbit'd2: is_wall <= 1'b1;
						`xbit'd3: is_wall <= 1'b1;
						`xbit'd4: is_wall <= 1'b1;
						`xbit'd5: is_wall <= 1'b1;
						`xbit'd6: is_wall <= 1'b1;
						`xbit'd7: is_wall <= 1'b1;
						`xbit'd8: is_wall <= 1'b1;
						`xbit'd9: is_wall <= 1'b1;
						`xbit'd10: is_wall <= 1'b1;
						`xbit'd11: is_wall <= 1'b1;
						`xbit'd12: is_wall <= 1'b1;
						`xbit'd13: is_wall <= 1'b1;
						`xbit'd14: is_wall <= 1'b1;
						`xbit'd15: is_wall <= 1'b1;
						`xbit'd16: is_wall <= 1'b1;
						`xbit'd17: is_wall <= 1'b1;
						`xbit'd18: is_wall <= 1'b1;
						`xbit'd19: is_wall <= 1'b1;
						`xbit'd20: is_wall <= 1'b1;
						`xbit'd21: is_wall <= 1'b1;
						`xbit'd22: is_wall <= 1'b1;
						`xbit'd23: is_wall <= 1'b1;
						`xbit'd24: is_wall <= 1'b1;
						`xbit'd25: is_wall <= 1'b1;
						`xbit'd26: is_wall <= 1'b1;
						`xbit'd27: is_wall <= 1'b1;
						`xbit'd28: is_wall <= 1'b1;
						`xbit'd29: is_wall <= 1'b1;
						`xbit'd30: is_wall <= 1'b1;
						`xbit'd31: is_wall <= 1'b1;
						`xbit'd32: is_wall <= 1'b1;
						`xbit'd33: is_wall <= 1'b1;
						`xbit'd34: is_wall <= 1'b1;
						`xbit'd35: is_wall <= 1'b1;
						`xbit'd36: is_wall <= 1'b1;
						`xbit'd37: is_wall <= 1'b1;
						`xbit'd38: is_wall <= 1'b1;
						`xbit'd39: is_wall <= 1'b1;
						`xbit'd40: is_wall <= 1'b1;
						`xbit'd41: is_wall <= 1'b1;
						`xbit'd42: is_wall <= 1'b1;
						`xbit'd43: is_wall <= 1'b1;
						`xbit'd44: is_wall <= 1'b1;
						`xbit'd45: is_wall <= 1'b1;
						`xbit'd46: is_wall <= 1'b1;
						`xbit'd47: is_wall <= 1'b1;
						`xbit'd48: is_wall <= 1'b1;
						`xbit'd49: is_wall <= 1'b1;
						`xbit'd50: is_wall <= 1'b1;
						`xbit'd51: is_wall <= 1'b1;
						`xbit'd52: is_wall <= 1'b1;
						`xbit'd53: is_wall <= 1'b1;
						`xbit'd54: is_wall <= 1'b1;
						`xbit'd55: is_wall <= 1'b1;
						`xbit'd56: is_wall <= 1'b1;
						`xbit'd57: is_wall <= 1'b1;
						`xbit'd58: is_wall <= 1'b1;
						`xbit'd59: is_wall <= 1'b1;
						`xbit'd60: is_wall <= 1'b1;
						`xbit'd61: is_wall <= 1'b1;
						`xbit'd62: is_wall <= 1'b1;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
				`ybit'd47: begin
					case(X)
						`xbit'd0: is_wall <= 1'b0;
						`xbit'd1: is_wall <= 1'b0;
						`xbit'd2: is_wall <= 1'b0;
						`xbit'd3: is_wall <= 1'b0;
						`xbit'd4: is_wall <= 1'b0;
						`xbit'd5: is_wall <= 1'b0;
						`xbit'd6: is_wall <= 1'b0;
						`xbit'd7: is_wall <= 1'b0;
						`xbit'd8: is_wall <= 1'b0;
						`xbit'd9: is_wall <= 1'b0;
						`xbit'd10: is_wall <= 1'b0;
						`xbit'd11: is_wall <= 1'b0;
						`xbit'd12: is_wall <= 1'b0;
						`xbit'd13: is_wall <= 1'b0;
						`xbit'd14: is_wall <= 1'b0;
						`xbit'd15: is_wall <= 1'b0;
						`xbit'd16: is_wall <= 1'b0;
						`xbit'd17: is_wall <= 1'b0;
						`xbit'd18: is_wall <= 1'b0;
						`xbit'd19: is_wall <= 1'b0;
						`xbit'd20: is_wall <= 1'b0;
						`xbit'd21: is_wall <= 1'b0;
						`xbit'd22: is_wall <= 1'b0;
						`xbit'd23: is_wall <= 1'b0;
						`xbit'd24: is_wall <= 1'b0;
						`xbit'd25: is_wall <= 1'b0;
						`xbit'd26: is_wall <= 1'b0;
						`xbit'd27: is_wall <= 1'b0;
						`xbit'd28: is_wall <= 1'b0;
						`xbit'd29: is_wall <= 1'b0;
						`xbit'd30: is_wall <= 1'b0;
						`xbit'd31: is_wall <= 1'b0;
						`xbit'd32: is_wall <= 1'b0;
						`xbit'd33: is_wall <= 1'b0;
						`xbit'd34: is_wall <= 1'b0;
						`xbit'd35: is_wall <= 1'b0;
						`xbit'd36: is_wall <= 1'b0;
						`xbit'd37: is_wall <= 1'b0;
						`xbit'd38: is_wall <= 1'b0;
						`xbit'd39: is_wall <= 1'b0;
						`xbit'd40: is_wall <= 1'b0;
						`xbit'd41: is_wall <= 1'b0;
						`xbit'd42: is_wall <= 1'b0;
						`xbit'd43: is_wall <= 1'b0;
						`xbit'd44: is_wall <= 1'b0;
						`xbit'd45: is_wall <= 1'b0;
						`xbit'd46: is_wall <= 1'b0;
						`xbit'd47: is_wall <= 1'b0;
						`xbit'd48: is_wall <= 1'b0;
						`xbit'd49: is_wall <= 1'b0;
						`xbit'd50: is_wall <= 1'b0;
						`xbit'd51: is_wall <= 1'b0;
						`xbit'd52: is_wall <= 1'b0;
						`xbit'd53: is_wall <= 1'b0;
						`xbit'd54: is_wall <= 1'b0;
						`xbit'd55: is_wall <= 1'b0;
						`xbit'd56: is_wall <= 1'b0;
						`xbit'd57: is_wall <= 1'b0;
						`xbit'd58: is_wall <= 1'b0;
						`xbit'd59: is_wall <= 1'b0;
						`xbit'd60: is_wall <= 1'b0;
						`xbit'd61: is_wall <= 1'b0;
						`xbit'd62: is_wall <= 1'b0;
						`xbit'd63: is_wall <= 1'b0;
					endcase
				end
			endcase
		end
	end

endmodule