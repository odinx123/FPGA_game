module filter(clk, rst, X, Y, data);

	parameter xbit = 10, ybit = 9;
	input clk, rst;
	input [xbit-1:0] X;
	input [ybit-1:0] Y;
	output data;
	reg data;

	wire [63:0] img[47:0];
	always@ (posedge clk, negedge rst) begin
		if (!rst) begin
			data <= 1'b0;
		end
		else begin
			if (img[Y][X] || img[Y-2][X] || img[Y+2]) begin
				data <= 1'b1;
			end
			else begin
				data <= 1'b0;
			end
		end
	end

	assign img[0][0] = 1'b0;
	assign img[0][1] = 1'b0;
	assign img[0][2] = 1'b0;
	assign img[0][3] = 1'b0;
	assign img[0][4] = 1'b0;
	assign img[0][5] = 1'b0;
	assign img[0][6] = 1'b0;
	assign img[0][7] = 1'b0;
	assign img[0][8] = 1'b0;
	assign img[0][9] = 1'b0;
	assign img[0][10] = 1'b0;
	assign img[0][11] = 1'b0;
	assign img[0][12] = 1'b0;
	assign img[0][13] = 1'b0;
	assign img[0][14] = 1'b0;
	assign img[0][15] = 1'b0;
	assign img[0][16] = 1'b0;
	assign img[0][17] = 1'b0;
	assign img[0][18] = 1'b0;
	assign img[0][19] = 1'b0;
	assign img[0][20] = 1'b0;
	assign img[0][21] = 1'b0;
	assign img[0][22] = 1'b0;
	assign img[0][23] = 1'b0;
	assign img[0][24] = 1'b0;
	assign img[0][25] = 1'b0;
	assign img[0][26] = 1'b0;
	assign img[0][27] = 1'b0;
	assign img[0][28] = 1'b0;
	assign img[0][29] = 1'b0;
	assign img[0][30] = 1'b0;
	assign img[0][31] = 1'b0;
	assign img[0][32] = 1'b0;
	assign img[0][33] = 1'b0;
	assign img[0][34] = 1'b0;
	assign img[0][35] = 1'b0;
	assign img[0][36] = 1'b0;
	assign img[0][37] = 1'b0;
	assign img[0][38] = 1'b0;
	assign img[0][39] = 1'b0;
	assign img[0][40] = 1'b0;
	assign img[0][41] = 1'b0;
	assign img[0][42] = 1'b0;
	assign img[0][43] = 1'b0;
	assign img[0][44] = 1'b0;
	assign img[0][45] = 1'b0;
	assign img[0][46] = 1'b0;
	assign img[0][47] = 1'b0;
	assign img[0][48] = 1'b0;
	assign img[0][49] = 1'b0;
	assign img[0][50] = 1'b0;
	assign img[0][51] = 1'b0;
	assign img[0][52] = 1'b0;
	assign img[0][53] = 1'b0;
	assign img[0][54] = 1'b0;
	assign img[0][55] = 1'b0;
	assign img[0][56] = 1'b0;
	assign img[0][57] = 1'b0;
	assign img[0][58] = 1'b0;
	assign img[0][59] = 1'b0;
	assign img[0][60] = 1'b0;
	assign img[0][61] = 1'b0;
	assign img[0][62] = 1'b0;
	assign img[0][63] = 1'b0;
	assign img[1][0] = 1'b0;
	assign img[1][1] = 1'b0;
	assign img[1][2] = 1'b0;
	assign img[1][3] = 1'b0;
	assign img[1][4] = 1'b0;
	assign img[1][5] = 1'b0;
	assign img[1][6] = 1'b0;
	assign img[1][7] = 1'b0;
	assign img[1][8] = 1'b0;
	assign img[1][9] = 1'b0;
	assign img[1][10] = 1'b0;
	assign img[1][11] = 1'b0;
	assign img[1][12] = 1'b0;
	assign img[1][13] = 1'b0;
	assign img[1][14] = 1'b0;
	assign img[1][15] = 1'b0;
	assign img[1][16] = 1'b0;
	assign img[1][17] = 1'b0;
	assign img[1][18] = 1'b0;
	assign img[1][19] = 1'b0;
	assign img[1][20] = 1'b0;
	assign img[1][21] = 1'b0;
	assign img[1][22] = 1'b0;
	assign img[1][23] = 1'b0;
	assign img[1][24] = 1'b0;
	assign img[1][25] = 1'b0;
	assign img[1][26] = 1'b0;
	assign img[1][27] = 1'b0;
	assign img[1][28] = 1'b0;
	assign img[1][29] = 1'b0;
	assign img[1][30] = 1'b0;
	assign img[1][31] = 1'b0;
	assign img[1][32] = 1'b0;
	assign img[1][33] = 1'b0;
	assign img[1][34] = 1'b0;
	assign img[1][35] = 1'b0;
	assign img[1][36] = 1'b0;
	assign img[1][37] = 1'b0;
	assign img[1][38] = 1'b0;
	assign img[1][39] = 1'b0;
	assign img[1][40] = 1'b0;
	assign img[1][41] = 1'b0;
	assign img[1][42] = 1'b0;
	assign img[1][43] = 1'b0;
	assign img[1][44] = 1'b0;
	assign img[1][45] = 1'b0;
	assign img[1][46] = 1'b0;
	assign img[1][47] = 1'b0;
	assign img[1][48] = 1'b0;
	assign img[1][49] = 1'b0;
	assign img[1][50] = 1'b0;
	assign img[1][51] = 1'b0;
	assign img[1][52] = 1'b0;
	assign img[1][53] = 1'b0;
	assign img[1][54] = 1'b0;
	assign img[1][55] = 1'b0;
	assign img[1][56] = 1'b0;
	assign img[1][57] = 1'b0;
	assign img[1][58] = 1'b0;
	assign img[1][59] = 1'b0;
	assign img[1][60] = 1'b0;
	assign img[1][61] = 1'b0;
	assign img[1][62] = 1'b0;
	assign img[1][63] = 1'b0;
	assign img[2][0] = 1'b0;
	assign img[2][1] = 1'b0;
	assign img[2][2] = 1'b0;
	assign img[2][3] = 1'b0;
	assign img[2][4] = 1'b0;
	assign img[2][5] = 1'b0;
	assign img[2][6] = 1'b0;
	assign img[2][7] = 1'b0;
	assign img[2][8] = 1'b0;
	assign img[2][9] = 1'b0;
	assign img[2][10] = 1'b0;
	assign img[2][11] = 1'b0;
	assign img[2][12] = 1'b0;
	assign img[2][13] = 1'b0;
	assign img[2][14] = 1'b0;
	assign img[2][15] = 1'b0;
	assign img[2][16] = 1'b0;
	assign img[2][17] = 1'b0;
	assign img[2][18] = 1'b0;
	assign img[2][19] = 1'b0;
	assign img[2][20] = 1'b0;
	assign img[2][21] = 1'b0;
	assign img[2][22] = 1'b0;
	assign img[2][23] = 1'b0;
	assign img[2][24] = 1'b0;
	assign img[2][25] = 1'b0;
	assign img[2][26] = 1'b0;
	assign img[2][27] = 1'b0;
	assign img[2][28] = 1'b0;
	assign img[2][29] = 1'b0;
	assign img[2][30] = 1'b0;
	assign img[2][31] = 1'b0;
	assign img[2][32] = 1'b0;
	assign img[2][33] = 1'b0;
	assign img[2][34] = 1'b0;
	assign img[2][35] = 1'b0;
	assign img[2][36] = 1'b0;
	assign img[2][37] = 1'b0;
	assign img[2][38] = 1'b0;
	assign img[2][39] = 1'b0;
	assign img[2][40] = 1'b0;
	assign img[2][41] = 1'b0;
	assign img[2][42] = 1'b0;
	assign img[2][43] = 1'b0;
	assign img[2][44] = 1'b0;
	assign img[2][45] = 1'b0;
	assign img[2][46] = 1'b0;
	assign img[2][47] = 1'b0;
	assign img[2][48] = 1'b0;
	assign img[2][49] = 1'b0;
	assign img[2][50] = 1'b0;
	assign img[2][51] = 1'b0;
	assign img[2][52] = 1'b0;
	assign img[2][53] = 1'b0;
	assign img[2][54] = 1'b0;
	assign img[2][55] = 1'b0;
	assign img[2][56] = 1'b0;
	assign img[2][57] = 1'b0;
	assign img[2][58] = 1'b0;
	assign img[2][59] = 1'b0;
	assign img[2][60] = 1'b0;
	assign img[2][61] = 1'b0;
	assign img[2][62] = 1'b0;
	assign img[2][63] = 1'b0;
	assign img[3][0] = 1'b0;
	assign img[3][1] = 1'b0;
	assign img[3][2] = 1'b0;
	assign img[3][3] = 1'b0;
	assign img[3][4] = 1'b0;
	assign img[3][5] = 1'b0;
	assign img[3][6] = 1'b0;
	assign img[3][7] = 1'b0;
	assign img[3][8] = 1'b0;
	assign img[3][9] = 1'b0;
	assign img[3][10] = 1'b0;
	assign img[3][11] = 1'b0;
	assign img[3][12] = 1'b0;
	assign img[3][13] = 1'b0;
	assign img[3][14] = 1'b0;
	assign img[3][15] = 1'b0;
	assign img[3][16] = 1'b0;
	assign img[3][17] = 1'b0;
	assign img[3][18] = 1'b0;
	assign img[3][19] = 1'b0;
	assign img[3][20] = 1'b0;
	assign img[3][21] = 1'b0;
	assign img[3][22] = 1'b0;
	assign img[3][23] = 1'b0;
	assign img[3][24] = 1'b0;
	assign img[3][25] = 1'b0;
	assign img[3][26] = 1'b0;
	assign img[3][27] = 1'b0;
	assign img[3][28] = 1'b0;
	assign img[3][29] = 1'b0;
	assign img[3][30] = 1'b0;
	assign img[3][31] = 1'b0;
	assign img[3][32] = 1'b0;
	assign img[3][33] = 1'b0;
	assign img[3][34] = 1'b0;
	assign img[3][35] = 1'b0;
	assign img[3][36] = 1'b0;
	assign img[3][37] = 1'b0;
	assign img[3][38] = 1'b0;
	assign img[3][39] = 1'b0;
	assign img[3][40] = 1'b0;
	assign img[3][41] = 1'b0;
	assign img[3][42] = 1'b0;
	assign img[3][43] = 1'b0;
	assign img[3][44] = 1'b0;
	assign img[3][45] = 1'b0;
	assign img[3][46] = 1'b0;
	assign img[3][47] = 1'b0;
	assign img[3][48] = 1'b0;
	assign img[3][49] = 1'b0;
	assign img[3][50] = 1'b0;
	assign img[3][51] = 1'b0;
	assign img[3][52] = 1'b0;
	assign img[3][53] = 1'b0;
	assign img[3][54] = 1'b0;
	assign img[3][55] = 1'b0;
	assign img[3][56] = 1'b0;
	assign img[3][57] = 1'b0;
	assign img[3][58] = 1'b0;
	assign img[3][59] = 1'b0;
	assign img[3][60] = 1'b0;
	assign img[3][61] = 1'b0;
	assign img[3][62] = 1'b0;
	assign img[3][63] = 1'b0;
	assign img[4][0] = 1'b0;
	assign img[4][1] = 1'b0;
	assign img[4][2] = 1'b0;
	assign img[4][3] = 1'b0;
	assign img[4][4] = 1'b0;
	assign img[4][5] = 1'b0;
	assign img[4][6] = 1'b0;
	assign img[4][7] = 1'b0;
	assign img[4][8] = 1'b0;
	assign img[4][9] = 1'b0;
	assign img[4][10] = 1'b0;
	assign img[4][11] = 1'b0;
	assign img[4][12] = 1'b0;
	assign img[4][13] = 1'b0;
	assign img[4][14] = 1'b0;
	assign img[4][15] = 1'b0;
	assign img[4][16] = 1'b0;
	assign img[4][17] = 1'b0;
	assign img[4][18] = 1'b0;
	assign img[4][19] = 1'b0;
	assign img[4][20] = 1'b0;
	assign img[4][21] = 1'b0;
	assign img[4][22] = 1'b0;
	assign img[4][23] = 1'b0;
	assign img[4][24] = 1'b0;
	assign img[4][25] = 1'b0;
	assign img[4][26] = 1'b0;
	assign img[4][27] = 1'b0;
	assign img[4][28] = 1'b0;
	assign img[4][29] = 1'b0;
	assign img[4][30] = 1'b0;
	assign img[4][31] = 1'b0;
	assign img[4][32] = 1'b0;
	assign img[4][33] = 1'b0;
	assign img[4][34] = 1'b0;
	assign img[4][35] = 1'b0;
	assign img[4][36] = 1'b0;
	assign img[4][37] = 1'b0;
	assign img[4][38] = 1'b0;
	assign img[4][39] = 1'b0;
	assign img[4][40] = 1'b0;
	assign img[4][41] = 1'b0;
	assign img[4][42] = 1'b0;
	assign img[4][43] = 1'b0;
	assign img[4][44] = 1'b0;
	assign img[4][45] = 1'b0;
	assign img[4][46] = 1'b0;
	assign img[4][47] = 1'b0;
	assign img[4][48] = 1'b0;
	assign img[4][49] = 1'b0;
	assign img[4][50] = 1'b0;
	assign img[4][51] = 1'b0;
	assign img[4][52] = 1'b0;
	assign img[4][53] = 1'b0;
	assign img[4][54] = 1'b0;
	assign img[4][55] = 1'b0;
	assign img[4][56] = 1'b0;
	assign img[4][57] = 1'b0;
	assign img[4][58] = 1'b0;
	assign img[4][59] = 1'b0;
	assign img[4][60] = 1'b0;
	assign img[4][61] = 1'b0;
	assign img[4][62] = 1'b0;
	assign img[4][63] = 1'b0;
	assign img[5][0] = 1'b0;
	assign img[5][1] = 1'b0;
	assign img[5][2] = 1'b0;
	assign img[5][3] = 1'b0;
	assign img[5][4] = 1'b0;
	assign img[5][5] = 1'b0;
	assign img[5][6] = 1'b0;
	assign img[5][7] = 1'b0;
	assign img[5][8] = 1'b0;
	assign img[5][9] = 1'b0;
	assign img[5][10] = 1'b0;
	assign img[5][11] = 1'b0;
	assign img[5][12] = 1'b0;
	assign img[5][13] = 1'b0;
	assign img[5][14] = 1'b0;
	assign img[5][15] = 1'b0;
	assign img[5][16] = 1'b0;
	assign img[5][17] = 1'b0;
	assign img[5][18] = 1'b0;
	assign img[5][19] = 1'b0;
	assign img[5][20] = 1'b0;
	assign img[5][21] = 1'b0;
	assign img[5][22] = 1'b0;
	assign img[5][23] = 1'b0;
	assign img[5][24] = 1'b0;
	assign img[5][25] = 1'b0;
	assign img[5][26] = 1'b0;
	assign img[5][27] = 1'b0;
	assign img[5][28] = 1'b0;
	assign img[5][29] = 1'b0;
	assign img[5][30] = 1'b0;
	assign img[5][31] = 1'b0;
	assign img[5][32] = 1'b0;
	assign img[5][33] = 1'b0;
	assign img[5][34] = 1'b0;
	assign img[5][35] = 1'b0;
	assign img[5][36] = 1'b0;
	assign img[5][37] = 1'b0;
	assign img[5][38] = 1'b0;
	assign img[5][39] = 1'b0;
	assign img[5][40] = 1'b0;
	assign img[5][41] = 1'b0;
	assign img[5][42] = 1'b0;
	assign img[5][43] = 1'b0;
	assign img[5][44] = 1'b0;
	assign img[5][45] = 1'b0;
	assign img[5][46] = 1'b0;
	assign img[5][47] = 1'b0;
	assign img[5][48] = 1'b0;
	assign img[5][49] = 1'b0;
	assign img[5][50] = 1'b0;
	assign img[5][51] = 1'b0;
	assign img[5][52] = 1'b0;
	assign img[5][53] = 1'b0;
	assign img[5][54] = 1'b0;
	assign img[5][55] = 1'b0;
	assign img[5][56] = 1'b0;
	assign img[5][57] = 1'b0;
	assign img[5][58] = 1'b0;
	assign img[5][59] = 1'b0;
	assign img[5][60] = 1'b0;
	assign img[5][61] = 1'b0;
	assign img[5][62] = 1'b0;
	assign img[5][63] = 1'b0;
	assign img[6][0] = 1'b0;
	assign img[6][1] = 1'b0;
	assign img[6][2] = 1'b0;
	assign img[6][3] = 1'b0;
	assign img[6][4] = 1'b0;
	assign img[6][5] = 1'b0;
	assign img[6][6] = 1'b0;
	assign img[6][7] = 1'b0;
	assign img[6][8] = 1'b0;
	assign img[6][9] = 1'b0;
	assign img[6][10] = 1'b0;
	assign img[6][11] = 1'b0;
	assign img[6][12] = 1'b0;
	assign img[6][13] = 1'b0;
	assign img[6][14] = 1'b0;
	assign img[6][15] = 1'b0;
	assign img[6][16] = 1'b0;
	assign img[6][17] = 1'b0;
	assign img[6][18] = 1'b0;
	assign img[6][19] = 1'b0;
	assign img[6][20] = 1'b0;
	assign img[6][21] = 1'b0;
	assign img[6][22] = 1'b0;
	assign img[6][23] = 1'b0;
	assign img[6][24] = 1'b0;
	assign img[6][25] = 1'b0;
	assign img[6][26] = 1'b0;
	assign img[6][27] = 1'b0;
	assign img[6][28] = 1'b0;
	assign img[6][29] = 1'b0;
	assign img[6][30] = 1'b0;
	assign img[6][31] = 1'b0;
	assign img[6][32] = 1'b0;
	assign img[6][33] = 1'b0;
	assign img[6][34] = 1'b0;
	assign img[6][35] = 1'b0;
	assign img[6][36] = 1'b0;
	assign img[6][37] = 1'b0;
	assign img[6][38] = 1'b0;
	assign img[6][39] = 1'b0;
	assign img[6][40] = 1'b0;
	assign img[6][41] = 1'b0;
	assign img[6][42] = 1'b0;
	assign img[6][43] = 1'b0;
	assign img[6][44] = 1'b0;
	assign img[6][45] = 1'b0;
	assign img[6][46] = 1'b0;
	assign img[6][47] = 1'b0;
	assign img[6][48] = 1'b0;
	assign img[6][49] = 1'b0;
	assign img[6][50] = 1'b0;
	assign img[6][51] = 1'b0;
	assign img[6][52] = 1'b0;
	assign img[6][53] = 1'b0;
	assign img[6][54] = 1'b0;
	assign img[6][55] = 1'b0;
	assign img[6][56] = 1'b0;
	assign img[6][57] = 1'b0;
	assign img[6][58] = 1'b0;
	assign img[6][59] = 1'b0;
	assign img[6][60] = 1'b0;
	assign img[6][61] = 1'b0;
	assign img[6][62] = 1'b0;
	assign img[6][63] = 1'b0;
	assign img[7][0] = 1'b0;
	assign img[7][1] = 1'b0;
	assign img[7][2] = 1'b0;
	assign img[7][3] = 1'b0;
	assign img[7][4] = 1'b0;
	assign img[7][5] = 1'b0;
	assign img[7][6] = 1'b0;
	assign img[7][7] = 1'b0;
	assign img[7][8] = 1'b0;
	assign img[7][9] = 1'b0;
	assign img[7][10] = 1'b0;
	assign img[7][11] = 1'b0;
	assign img[7][12] = 1'b0;
	assign img[7][13] = 1'b0;
	assign img[7][14] = 1'b0;
	assign img[7][15] = 1'b0;
	assign img[7][16] = 1'b0;
	assign img[7][17] = 1'b0;
	assign img[7][18] = 1'b0;
	assign img[7][19] = 1'b0;
	assign img[7][20] = 1'b0;
	assign img[7][21] = 1'b0;
	assign img[7][22] = 1'b0;
	assign img[7][23] = 1'b0;
	assign img[7][24] = 1'b0;
	assign img[7][25] = 1'b0;
	assign img[7][26] = 1'b0;
	assign img[7][27] = 1'b0;
	assign img[7][28] = 1'b0;
	assign img[7][29] = 1'b0;
	assign img[7][30] = 1'b0;
	assign img[7][31] = 1'b0;
	assign img[7][32] = 1'b0;
	assign img[7][33] = 1'b0;
	assign img[7][34] = 1'b0;
	assign img[7][35] = 1'b0;
	assign img[7][36] = 1'b0;
	assign img[7][37] = 1'b0;
	assign img[7][38] = 1'b0;
	assign img[7][39] = 1'b0;
	assign img[7][40] = 1'b0;
	assign img[7][41] = 1'b0;
	assign img[7][42] = 1'b0;
	assign img[7][43] = 1'b0;
	assign img[7][44] = 1'b0;
	assign img[7][45] = 1'b0;
	assign img[7][46] = 1'b0;
	assign img[7][47] = 1'b0;
	assign img[7][48] = 1'b0;
	assign img[7][49] = 1'b0;
	assign img[7][50] = 1'b0;
	assign img[7][51] = 1'b0;
	assign img[7][52] = 1'b0;
	assign img[7][53] = 1'b0;
	assign img[7][54] = 1'b0;
	assign img[7][55] = 1'b0;
	assign img[7][56] = 1'b0;
	assign img[7][57] = 1'b0;
	assign img[7][58] = 1'b0;
	assign img[7][59] = 1'b0;
	assign img[7][60] = 1'b0;
	assign img[7][61] = 1'b0;
	assign img[7][62] = 1'b0;
	assign img[7][63] = 1'b0;
	assign img[8][0] = 1'b0;
	assign img[8][1] = 1'b0;
	assign img[8][2] = 1'b0;
	assign img[8][3] = 1'b0;
	assign img[8][4] = 1'b0;
	assign img[8][5] = 1'b0;
	assign img[8][6] = 1'b0;
	assign img[8][7] = 1'b0;
	assign img[8][8] = 1'b0;
	assign img[8][9] = 1'b0;
	assign img[8][10] = 1'b0;
	assign img[8][11] = 1'b0;
	assign img[8][12] = 1'b0;
	assign img[8][13] = 1'b0;
	assign img[8][14] = 1'b0;
	assign img[8][15] = 1'b0;
	assign img[8][16] = 1'b0;
	assign img[8][17] = 1'b0;
	assign img[8][18] = 1'b0;
	assign img[8][19] = 1'b0;
	assign img[8][20] = 1'b0;
	assign img[8][21] = 1'b0;
	assign img[8][22] = 1'b0;
	assign img[8][23] = 1'b0;
	assign img[8][24] = 1'b0;
	assign img[8][25] = 1'b0;
	assign img[8][26] = 1'b0;
	assign img[8][27] = 1'b0;
	assign img[8][28] = 1'b0;
	assign img[8][29] = 1'b0;
	assign img[8][30] = 1'b0;
	assign img[8][31] = 1'b0;
	assign img[8][32] = 1'b0;
	assign img[8][33] = 1'b0;
	assign img[8][34] = 1'b0;
	assign img[8][35] = 1'b0;
	assign img[8][36] = 1'b0;
	assign img[8][37] = 1'b0;
	assign img[8][38] = 1'b0;
	assign img[8][39] = 1'b0;
	assign img[8][40] = 1'b0;
	assign img[8][41] = 1'b0;
	assign img[8][42] = 1'b0;
	assign img[8][43] = 1'b0;
	assign img[8][44] = 1'b0;
	assign img[8][45] = 1'b0;
	assign img[8][46] = 1'b0;
	assign img[8][47] = 1'b0;
	assign img[8][48] = 1'b0;
	assign img[8][49] = 1'b0;
	assign img[8][50] = 1'b0;
	assign img[8][51] = 1'b0;
	assign img[8][52] = 1'b0;
	assign img[8][53] = 1'b0;
	assign img[8][54] = 1'b0;
	assign img[8][55] = 1'b0;
	assign img[8][56] = 1'b0;
	assign img[8][57] = 1'b0;
	assign img[8][58] = 1'b0;
	assign img[8][59] = 1'b0;
	assign img[8][60] = 1'b0;
	assign img[8][61] = 1'b0;
	assign img[8][62] = 1'b0;
	assign img[8][63] = 1'b0;
	assign img[9][0] = 1'b0;
	assign img[9][1] = 1'b0;
	assign img[9][2] = 1'b0;
	assign img[9][3] = 1'b0;
	assign img[9][4] = 1'b0;
	assign img[9][5] = 1'b0;
	assign img[9][6] = 1'b0;
	assign img[9][7] = 1'b0;
	assign img[9][8] = 1'b0;
	assign img[9][9] = 1'b0;
	assign img[9][10] = 1'b0;
	assign img[9][11] = 1'b0;
	assign img[9][12] = 1'b0;
	assign img[9][13] = 1'b0;
	assign img[9][14] = 1'b0;
	assign img[9][15] = 1'b0;
	assign img[9][16] = 1'b0;
	assign img[9][17] = 1'b0;
	assign img[9][18] = 1'b0;
	assign img[9][19] = 1'b0;
	assign img[9][20] = 1'b0;
	assign img[9][21] = 1'b0;
	assign img[9][22] = 1'b0;
	assign img[9][23] = 1'b0;
	assign img[9][24] = 1'b0;
	assign img[9][25] = 1'b0;
	assign img[9][26] = 1'b0;
	assign img[9][27] = 1'b0;
	assign img[9][28] = 1'b0;
	assign img[9][29] = 1'b0;
	assign img[9][30] = 1'b0;
	assign img[9][31] = 1'b0;
	assign img[9][32] = 1'b0;
	assign img[9][33] = 1'b0;
	assign img[9][34] = 1'b0;
	assign img[9][35] = 1'b0;
	assign img[9][36] = 1'b0;
	assign img[9][37] = 1'b0;
	assign img[9][38] = 1'b0;
	assign img[9][39] = 1'b0;
	assign img[9][40] = 1'b0;
	assign img[9][41] = 1'b0;
	assign img[9][42] = 1'b0;
	assign img[9][43] = 1'b0;
	assign img[9][44] = 1'b0;
	assign img[9][45] = 1'b0;
	assign img[9][46] = 1'b0;
	assign img[9][47] = 1'b0;
	assign img[9][48] = 1'b0;
	assign img[9][49] = 1'b0;
	assign img[9][50] = 1'b0;
	assign img[9][51] = 1'b0;
	assign img[9][52] = 1'b0;
	assign img[9][53] = 1'b0;
	assign img[9][54] = 1'b0;
	assign img[9][55] = 1'b0;
	assign img[9][56] = 1'b0;
	assign img[9][57] = 1'b0;
	assign img[9][58] = 1'b0;
	assign img[9][59] = 1'b0;
	assign img[9][60] = 1'b0;
	assign img[9][61] = 1'b0;
	assign img[9][62] = 1'b0;
	assign img[9][63] = 1'b0;
	assign img[10][0] = 1'b0;
	assign img[10][1] = 1'b0;
	assign img[10][2] = 1'b0;
	assign img[10][3] = 1'b0;
	assign img[10][4] = 1'b0;
	assign img[10][5] = 1'b0;
	assign img[10][6] = 1'b0;
	assign img[10][7] = 1'b0;
	assign img[10][8] = 1'b0;
	assign img[10][9] = 1'b0;
	assign img[10][10] = 1'b0;
	assign img[10][11] = 1'b0;
	assign img[10][12] = 1'b0;
	assign img[10][13] = 1'b0;
	assign img[10][14] = 1'b0;
	assign img[10][15] = 1'b0;
	assign img[10][16] = 1'b0;
	assign img[10][17] = 1'b0;
	assign img[10][18] = 1'b0;
	assign img[10][19] = 1'b0;
	assign img[10][20] = 1'b0;
	assign img[10][21] = 1'b0;
	assign img[10][22] = 1'b0;
	assign img[10][23] = 1'b0;
	assign img[10][24] = 1'b0;
	assign img[10][25] = 1'b0;
	assign img[10][26] = 1'b0;
	assign img[10][27] = 1'b0;
	assign img[10][28] = 1'b0;
	assign img[10][29] = 1'b0;
	assign img[10][30] = 1'b0;
	assign img[10][31] = 1'b0;
	assign img[10][32] = 1'b0;
	assign img[10][33] = 1'b0;
	assign img[10][34] = 1'b0;
	assign img[10][35] = 1'b0;
	assign img[10][36] = 1'b0;
	assign img[10][37] = 1'b0;
	assign img[10][38] = 1'b0;
	assign img[10][39] = 1'b0;
	assign img[10][40] = 1'b0;
	assign img[10][41] = 1'b0;
	assign img[10][42] = 1'b0;
	assign img[10][43] = 1'b0;
	assign img[10][44] = 1'b0;
	assign img[10][45] = 1'b0;
	assign img[10][46] = 1'b0;
	assign img[10][47] = 1'b0;
	assign img[10][48] = 1'b0;
	assign img[10][49] = 1'b0;
	assign img[10][50] = 1'b0;
	assign img[10][51] = 1'b0;
	assign img[10][52] = 1'b1;
	assign img[10][53] = 1'b0;
	assign img[10][54] = 1'b0;
	assign img[10][55] = 1'b0;
	assign img[10][56] = 1'b0;
	assign img[10][57] = 1'b0;
	assign img[10][58] = 1'b0;
	assign img[10][59] = 1'b0;
	assign img[10][60] = 1'b0;
	assign img[10][61] = 1'b0;
	assign img[10][62] = 1'b0;
	assign img[10][63] = 1'b0;
	assign img[11][0] = 1'b0;
	assign img[11][1] = 1'b0;
	assign img[11][2] = 1'b0;
	assign img[11][3] = 1'b0;
	assign img[11][4] = 1'b0;
	assign img[11][5] = 1'b0;
	assign img[11][6] = 1'b0;
	assign img[11][7] = 1'b0;
	assign img[11][8] = 1'b0;
	assign img[11][9] = 1'b1;
	assign img[11][10] = 1'b0;
	assign img[11][11] = 1'b0;
	assign img[11][12] = 1'b0;
	assign img[11][13] = 1'b0;
	assign img[11][14] = 1'b0;
	assign img[11][15] = 1'b0;
	assign img[11][16] = 1'b0;
	assign img[11][17] = 1'b0;
	assign img[11][18] = 1'b0;
	assign img[11][19] = 1'b0;
	assign img[11][20] = 1'b0;
	assign img[11][21] = 1'b0;
	assign img[11][22] = 1'b0;
	assign img[11][23] = 1'b0;
	assign img[11][24] = 1'b0;
	assign img[11][25] = 1'b0;
	assign img[11][26] = 1'b0;
	assign img[11][27] = 1'b0;
	assign img[11][28] = 1'b0;
	assign img[11][29] = 1'b0;
	assign img[11][30] = 1'b0;
	assign img[11][31] = 1'b0;
	assign img[11][32] = 1'b0;
	assign img[11][33] = 1'b0;
	assign img[11][34] = 1'b0;
	assign img[11][35] = 1'b0;
	assign img[11][36] = 1'b0;
	assign img[11][37] = 1'b0;
	assign img[11][38] = 1'b0;
	assign img[11][39] = 1'b0;
	assign img[11][40] = 1'b0;
	assign img[11][41] = 1'b0;
	assign img[11][42] = 1'b0;
	assign img[11][43] = 1'b0;
	assign img[11][44] = 1'b0;
	assign img[11][45] = 1'b0;
	assign img[11][46] = 1'b0;
	assign img[11][47] = 1'b0;
	assign img[11][48] = 1'b0;
	assign img[11][49] = 1'b0;
	assign img[11][50] = 1'b0;
	assign img[11][51] = 1'b0;
	assign img[11][52] = 1'b0;
	assign img[11][53] = 1'b0;
	assign img[11][54] = 1'b0;
	assign img[11][55] = 1'b0;
	assign img[11][56] = 1'b0;
	assign img[11][57] = 1'b0;
	assign img[11][58] = 1'b0;
	assign img[11][59] = 1'b0;
	assign img[11][60] = 1'b0;
	assign img[11][61] = 1'b0;
	assign img[11][62] = 1'b0;
	assign img[11][63] = 1'b0;
	assign img[12][0] = 1'b0;
	assign img[12][1] = 1'b0;
	assign img[12][2] = 1'b0;
	assign img[12][3] = 1'b0;
	assign img[12][4] = 1'b0;
	assign img[12][5] = 1'b0;
	assign img[12][6] = 1'b0;
	assign img[12][7] = 1'b0;
	assign img[12][8] = 1'b0;
	assign img[12][9] = 1'b0;
	assign img[12][10] = 1'b0;
	assign img[12][11] = 1'b0;
	assign img[12][12] = 1'b0;
	assign img[12][13] = 1'b0;
	assign img[12][14] = 1'b0;
	assign img[12][15] = 1'b0;
	assign img[12][16] = 1'b0;
	assign img[12][17] = 1'b0;
	assign img[12][18] = 1'b0;
	assign img[12][19] = 1'b0;
	assign img[12][20] = 1'b0;
	assign img[12][21] = 1'b0;
	assign img[12][22] = 1'b0;
	assign img[12][23] = 1'b0;
	assign img[12][24] = 1'b0;
	assign img[12][25] = 1'b0;
	assign img[12][26] = 1'b0;
	assign img[12][27] = 1'b0;
	assign img[12][28] = 1'b0;
	assign img[12][29] = 1'b0;
	assign img[12][30] = 1'b0;
	assign img[12][31] = 1'b0;
	assign img[12][32] = 1'b0;
	assign img[12][33] = 1'b0;
	assign img[12][34] = 1'b0;
	assign img[12][35] = 1'b0;
	assign img[12][36] = 1'b0;
	assign img[12][37] = 1'b0;
	assign img[12][38] = 1'b0;
	assign img[12][39] = 1'b0;
	assign img[12][40] = 1'b0;
	assign img[12][41] = 1'b0;
	assign img[12][42] = 1'b0;
	assign img[12][43] = 1'b0;
	assign img[12][44] = 1'b0;
	assign img[12][45] = 1'b0;
	assign img[12][46] = 1'b0;
	assign img[12][47] = 1'b0;
	assign img[12][48] = 1'b0;
	assign img[12][49] = 1'b0;
	assign img[12][50] = 1'b0;
	assign img[12][51] = 1'b0;
	assign img[12][52] = 1'b0;
	assign img[12][53] = 1'b0;
	assign img[12][54] = 1'b0;
	assign img[12][55] = 1'b0;
	assign img[12][56] = 1'b0;
	assign img[12][57] = 1'b0;
	assign img[12][58] = 1'b0;
	assign img[12][59] = 1'b0;
	assign img[12][60] = 1'b0;
	assign img[12][61] = 1'b0;
	assign img[12][62] = 1'b0;
	assign img[12][63] = 1'b0;
	assign img[13][0] = 1'b0;
	assign img[13][1] = 1'b0;
	assign img[13][2] = 1'b0;
	assign img[13][3] = 1'b0;
	assign img[13][4] = 1'b0;
	assign img[13][5] = 1'b0;
	assign img[13][6] = 1'b0;
	assign img[13][7] = 1'b0;
	assign img[13][8] = 1'b0;
	assign img[13][9] = 1'b0;
	assign img[13][10] = 1'b0;
	assign img[13][11] = 1'b0;
	assign img[13][12] = 1'b0;
	assign img[13][13] = 1'b0;
	assign img[13][14] = 1'b0;
	assign img[13][15] = 1'b0;
	assign img[13][16] = 1'b0;
	assign img[13][17] = 1'b0;
	assign img[13][18] = 1'b0;
	assign img[13][19] = 1'b0;
	assign img[13][20] = 1'b0;
	assign img[13][21] = 1'b0;
	assign img[13][22] = 1'b0;
	assign img[13][23] = 1'b0;
	assign img[13][24] = 1'b0;
	assign img[13][25] = 1'b0;
	assign img[13][26] = 1'b0;
	assign img[13][27] = 1'b0;
	assign img[13][28] = 1'b0;
	assign img[13][29] = 1'b0;
	assign img[13][30] = 1'b0;
	assign img[13][31] = 1'b0;
	assign img[13][32] = 1'b0;
	assign img[13][33] = 1'b0;
	assign img[13][34] = 1'b0;
	assign img[13][35] = 1'b0;
	assign img[13][36] = 1'b0;
	assign img[13][37] = 1'b0;
	assign img[13][38] = 1'b0;
	assign img[13][39] = 1'b0;
	assign img[13][40] = 1'b0;
	assign img[13][41] = 1'b0;
	assign img[13][42] = 1'b0;
	assign img[13][43] = 1'b0;
	assign img[13][44] = 1'b0;
	assign img[13][45] = 1'b0;
	assign img[13][46] = 1'b0;
	assign img[13][47] = 1'b0;
	assign img[13][48] = 1'b0;
	assign img[13][49] = 1'b0;
	assign img[13][50] = 1'b0;
	assign img[13][51] = 1'b0;
	assign img[13][52] = 1'b0;
	assign img[13][53] = 1'b0;
	assign img[13][54] = 1'b0;
	assign img[13][55] = 1'b0;
	assign img[13][56] = 1'b0;
	assign img[13][57] = 1'b0;
	assign img[13][58] = 1'b0;
	assign img[13][59] = 1'b0;
	assign img[13][60] = 1'b0;
	assign img[13][61] = 1'b0;
	assign img[13][62] = 1'b0;
	assign img[13][63] = 1'b0;
	assign img[14][0] = 1'b0;
	assign img[14][1] = 1'b0;
	assign img[14][2] = 1'b0;
	assign img[14][3] = 1'b0;
	assign img[14][4] = 1'b0;
	assign img[14][5] = 1'b0;
	assign img[14][6] = 1'b0;
	assign img[14][7] = 1'b0;
	assign img[14][8] = 1'b0;
	assign img[14][9] = 1'b0;
	assign img[14][10] = 1'b0;
	assign img[14][11] = 1'b0;
	assign img[14][12] = 1'b0;
	assign img[14][13] = 1'b0;
	assign img[14][14] = 1'b0;
	assign img[14][15] = 1'b0;
	assign img[14][16] = 1'b0;
	assign img[14][17] = 1'b0;
	assign img[14][18] = 1'b0;
	assign img[14][19] = 1'b0;
	assign img[14][20] = 1'b0;
	assign img[14][21] = 1'b0;
	assign img[14][22] = 1'b0;
	assign img[14][23] = 1'b0;
	assign img[14][24] = 1'b0;
	assign img[14][25] = 1'b0;
	assign img[14][26] = 1'b0;
	assign img[14][27] = 1'b0;
	assign img[14][28] = 1'b0;
	assign img[14][29] = 1'b0;
	assign img[14][30] = 1'b0;
	assign img[14][31] = 1'b0;
	assign img[14][32] = 1'b0;
	assign img[14][33] = 1'b0;
	assign img[14][34] = 1'b0;
	assign img[14][35] = 1'b0;
	assign img[14][36] = 1'b0;
	assign img[14][37] = 1'b0;
	assign img[14][38] = 1'b0;
	assign img[14][39] = 1'b0;
	assign img[14][40] = 1'b0;
	assign img[14][41] = 1'b0;
	assign img[14][42] = 1'b0;
	assign img[14][43] = 1'b0;
	assign img[14][44] = 1'b0;
	assign img[14][45] = 1'b0;
	assign img[14][46] = 1'b0;
	assign img[14][47] = 1'b0;
	assign img[14][48] = 1'b0;
	assign img[14][49] = 1'b0;
	assign img[14][50] = 1'b0;
	assign img[14][51] = 1'b0;
	assign img[14][52] = 1'b0;
	assign img[14][53] = 1'b0;
	assign img[14][54] = 1'b0;
	assign img[14][55] = 1'b0;
	assign img[14][56] = 1'b0;
	assign img[14][57] = 1'b0;
	assign img[14][58] = 1'b0;
	assign img[14][59] = 1'b0;
	assign img[14][60] = 1'b0;
	assign img[14][61] = 1'b0;
	assign img[14][62] = 1'b0;
	assign img[14][63] = 1'b0;
	assign img[15][0] = 1'b0;
	assign img[15][1] = 1'b0;
	assign img[15][2] = 1'b0;
	assign img[15][3] = 1'b0;
	assign img[15][4] = 1'b0;
	assign img[15][5] = 1'b0;
	assign img[15][6] = 1'b0;
	assign img[15][7] = 1'b0;
	assign img[15][8] = 1'b0;
	assign img[15][9] = 1'b0;
	assign img[15][10] = 1'b0;
	assign img[15][11] = 1'b0;
	assign img[15][12] = 1'b0;
	assign img[15][13] = 1'b0;
	assign img[15][14] = 1'b0;
	assign img[15][15] = 1'b0;
	assign img[15][16] = 1'b0;
	assign img[15][17] = 1'b0;
	assign img[15][18] = 1'b0;
	assign img[15][19] = 1'b0;
	assign img[15][20] = 1'b0;
	assign img[15][21] = 1'b0;
	assign img[15][22] = 1'b0;
	assign img[15][23] = 1'b0;
	assign img[15][24] = 1'b0;
	assign img[15][25] = 1'b0;
	assign img[15][26] = 1'b0;
	assign img[15][27] = 1'b0;
	assign img[15][28] = 1'b0;
	assign img[15][29] = 1'b0;
	assign img[15][30] = 1'b0;
	assign img[15][31] = 1'b0;
	assign img[15][32] = 1'b0;
	assign img[15][33] = 1'b0;
	assign img[15][34] = 1'b0;
	assign img[15][35] = 1'b0;
	assign img[15][36] = 1'b0;
	assign img[15][37] = 1'b0;
	assign img[15][38] = 1'b0;
	assign img[15][39] = 1'b0;
	assign img[15][40] = 1'b0;
	assign img[15][41] = 1'b0;
	assign img[15][42] = 1'b0;
	assign img[15][43] = 1'b0;
	assign img[15][44] = 1'b0;
	assign img[15][45] = 1'b0;
	assign img[15][46] = 1'b0;
	assign img[15][47] = 1'b0;
	assign img[15][48] = 1'b0;
	assign img[15][49] = 1'b0;
	assign img[15][50] = 1'b0;
	assign img[15][51] = 1'b0;
	assign img[15][52] = 1'b0;
	assign img[15][53] = 1'b0;
	assign img[15][54] = 1'b0;
	assign img[15][55] = 1'b0;
	assign img[15][56] = 1'b0;
	assign img[15][57] = 1'b0;
	assign img[15][58] = 1'b0;
	assign img[15][59] = 1'b0;
	assign img[15][60] = 1'b0;
	assign img[15][61] = 1'b0;
	assign img[15][62] = 1'b1;
	assign img[15][63] = 1'b0;
	assign img[16][0] = 1'b0;
	assign img[16][1] = 1'b0;
	assign img[16][2] = 1'b0;
	assign img[16][3] = 1'b0;
	assign img[16][4] = 1'b0;
	assign img[16][5] = 1'b0;
	assign img[16][6] = 1'b0;
	assign img[16][7] = 1'b0;
	assign img[16][8] = 1'b0;
	assign img[16][9] = 1'b0;
	assign img[16][10] = 1'b0;
	assign img[16][11] = 1'b0;
	assign img[16][12] = 1'b0;
	assign img[16][13] = 1'b0;
	assign img[16][14] = 1'b0;
	assign img[16][15] = 1'b0;
	assign img[16][16] = 1'b0;
	assign img[16][17] = 1'b0;
	assign img[16][18] = 1'b0;
	assign img[16][19] = 1'b0;
	assign img[16][20] = 1'b0;
	assign img[16][21] = 1'b0;
	assign img[16][22] = 1'b0;
	assign img[16][23] = 1'b0;
	assign img[16][24] = 1'b0;
	assign img[16][25] = 1'b0;
	assign img[16][26] = 1'b0;
	assign img[16][27] = 1'b0;
	assign img[16][28] = 1'b0;
	assign img[16][29] = 1'b0;
	assign img[16][30] = 1'b0;
	assign img[16][31] = 1'b0;
	assign img[16][32] = 1'b0;
	assign img[16][33] = 1'b0;
	assign img[16][34] = 1'b0;
	assign img[16][35] = 1'b0;
	assign img[16][36] = 1'b0;
	assign img[16][37] = 1'b0;
	assign img[16][38] = 1'b0;
	assign img[16][39] = 1'b0;
	assign img[16][40] = 1'b0;
	assign img[16][41] = 1'b0;
	assign img[16][42] = 1'b0;
	assign img[16][43] = 1'b0;
	assign img[16][44] = 1'b0;
	assign img[16][45] = 1'b0;
	assign img[16][46] = 1'b0;
	assign img[16][47] = 1'b0;
	assign img[16][48] = 1'b0;
	assign img[16][49] = 1'b0;
	assign img[16][50] = 1'b0;
	assign img[16][51] = 1'b0;
	assign img[16][52] = 1'b0;
	assign img[16][53] = 1'b0;
	assign img[16][54] = 1'b0;
	assign img[16][55] = 1'b0;
	assign img[16][56] = 1'b0;
	assign img[16][57] = 1'b0;
	assign img[16][58] = 1'b0;
	assign img[16][59] = 1'b0;
	assign img[16][60] = 1'b0;
	assign img[16][61] = 1'b0;
	assign img[16][62] = 1'b0;
	assign img[16][63] = 1'b0;
	assign img[17][0] = 1'b0;
	assign img[17][1] = 1'b0;
	assign img[17][2] = 1'b0;
	assign img[17][3] = 1'b0;
	assign img[17][4] = 1'b0;
	assign img[17][5] = 1'b0;
	assign img[17][6] = 1'b0;
	assign img[17][7] = 1'b0;
	assign img[17][8] = 1'b0;
	assign img[17][9] = 1'b0;
	assign img[17][10] = 1'b0;
	assign img[17][11] = 1'b0;
	assign img[17][12] = 1'b0;
	assign img[17][13] = 1'b0;
	assign img[17][14] = 1'b0;
	assign img[17][15] = 1'b0;
	assign img[17][16] = 1'b0;
	assign img[17][17] = 1'b0;
	assign img[17][18] = 1'b0;
	assign img[17][19] = 1'b0;
	assign img[17][20] = 1'b0;
	assign img[17][21] = 1'b0;
	assign img[17][22] = 1'b0;
	assign img[17][23] = 1'b0;
	assign img[17][24] = 1'b0;
	assign img[17][25] = 1'b0;
	assign img[17][26] = 1'b0;
	assign img[17][27] = 1'b0;
	assign img[17][28] = 1'b0;
	assign img[17][29] = 1'b0;
	assign img[17][30] = 1'b0;
	assign img[17][31] = 1'b0;
	assign img[17][32] = 1'b0;
	assign img[17][33] = 1'b0;
	assign img[17][34] = 1'b0;
	assign img[17][35] = 1'b0;
	assign img[17][36] = 1'b0;
	assign img[17][37] = 1'b0;
	assign img[17][38] = 1'b0;
	assign img[17][39] = 1'b0;
	assign img[17][40] = 1'b0;
	assign img[17][41] = 1'b0;
	assign img[17][42] = 1'b0;
	assign img[17][43] = 1'b0;
	assign img[17][44] = 1'b0;
	assign img[17][45] = 1'b0;
	assign img[17][46] = 1'b0;
	assign img[17][47] = 1'b0;
	assign img[17][48] = 1'b0;
	assign img[17][49] = 1'b0;
	assign img[17][50] = 1'b0;
	assign img[17][51] = 1'b0;
	assign img[17][52] = 1'b0;
	assign img[17][53] = 1'b0;
	assign img[17][54] = 1'b0;
	assign img[17][55] = 1'b0;
	assign img[17][56] = 1'b0;
	assign img[17][57] = 1'b0;
	assign img[17][58] = 1'b0;
	assign img[17][59] = 1'b0;
	assign img[17][60] = 1'b0;
	assign img[17][61] = 1'b0;
	assign img[17][62] = 1'b0;
	assign img[17][63] = 1'b0;
	assign img[18][0] = 1'b0;
	assign img[18][1] = 1'b0;
	assign img[18][2] = 1'b0;
	assign img[18][3] = 1'b0;
	assign img[18][4] = 1'b0;
	assign img[18][5] = 1'b0;
	assign img[18][6] = 1'b0;
	assign img[18][7] = 1'b0;
	assign img[18][8] = 1'b0;
	assign img[18][9] = 1'b0;
	assign img[18][10] = 1'b0;
	assign img[18][11] = 1'b0;
	assign img[18][12] = 1'b0;
	assign img[18][13] = 1'b0;
	assign img[18][14] = 1'b0;
	assign img[18][15] = 1'b0;
	assign img[18][16] = 1'b0;
	assign img[18][17] = 1'b1;
	assign img[18][18] = 1'b0;
	assign img[18][19] = 1'b0;
	assign img[18][20] = 1'b0;
	assign img[18][21] = 1'b0;
	assign img[18][22] = 1'b0;
	assign img[18][23] = 1'b0;
	assign img[18][24] = 1'b0;
	assign img[18][25] = 1'b0;
	assign img[18][26] = 1'b0;
	assign img[18][27] = 1'b0;
	assign img[18][28] = 1'b0;
	assign img[18][29] = 1'b0;
	assign img[18][30] = 1'b0;
	assign img[18][31] = 1'b0;
	assign img[18][32] = 1'b0;
	assign img[18][33] = 1'b0;
	assign img[18][34] = 1'b0;
	assign img[18][35] = 1'b0;
	assign img[18][36] = 1'b0;
	assign img[18][37] = 1'b0;
	assign img[18][38] = 1'b0;
	assign img[18][39] = 1'b0;
	assign img[18][40] = 1'b0;
	assign img[18][41] = 1'b0;
	assign img[18][42] = 1'b0;
	assign img[18][43] = 1'b0;
	assign img[18][44] = 1'b0;
	assign img[18][45] = 1'b0;
	assign img[18][46] = 1'b0;
	assign img[18][47] = 1'b0;
	assign img[18][48] = 1'b0;
	assign img[18][49] = 1'b0;
	assign img[18][50] = 1'b0;
	assign img[18][51] = 1'b0;
	assign img[18][52] = 1'b0;
	assign img[18][53] = 1'b0;
	assign img[18][54] = 1'b0;
	assign img[18][55] = 1'b0;
	assign img[18][56] = 1'b0;
	assign img[18][57] = 1'b0;
	assign img[18][58] = 1'b0;
	assign img[18][59] = 1'b0;
	assign img[18][60] = 1'b0;
	assign img[18][61] = 1'b0;
	assign img[18][62] = 1'b0;
	assign img[18][63] = 1'b0;
	assign img[19][0] = 1'b0;
	assign img[19][1] = 1'b0;
	assign img[19][2] = 1'b0;
	assign img[19][3] = 1'b0;
	assign img[19][4] = 1'b0;
	assign img[19][5] = 1'b0;
	assign img[19][6] = 1'b0;
	assign img[19][7] = 1'b0;
	assign img[19][8] = 1'b0;
	assign img[19][9] = 1'b0;
	assign img[19][10] = 1'b0;
	assign img[19][11] = 1'b0;
	assign img[19][12] = 1'b0;
	assign img[19][13] = 1'b1;
	assign img[19][14] = 1'b0;
	assign img[19][15] = 1'b0;
	assign img[19][16] = 1'b0;
	assign img[19][17] = 1'b0;
	assign img[19][18] = 1'b0;
	assign img[19][19] = 1'b0;
	assign img[19][20] = 1'b0;
	assign img[19][21] = 1'b0;
	assign img[19][22] = 1'b0;
	assign img[19][23] = 1'b0;
	assign img[19][24] = 1'b0;
	assign img[19][25] = 1'b0;
	assign img[19][26] = 1'b0;
	assign img[19][27] = 1'b0;
	assign img[19][28] = 1'b0;
	assign img[19][29] = 1'b0;
	assign img[19][30] = 1'b0;
	assign img[19][31] = 1'b0;
	assign img[19][32] = 1'b0;
	assign img[19][33] = 1'b0;
	assign img[19][34] = 1'b0;
	assign img[19][35] = 1'b0;
	assign img[19][36] = 1'b0;
	assign img[19][37] = 1'b0;
	assign img[19][38] = 1'b0;
	assign img[19][39] = 1'b0;
	assign img[19][40] = 1'b0;
	assign img[19][41] = 1'b0;
	assign img[19][42] = 1'b0;
	assign img[19][43] = 1'b0;
	assign img[19][44] = 1'b0;
	assign img[19][45] = 1'b0;
	assign img[19][46] = 1'b0;
	assign img[19][47] = 1'b0;
	assign img[19][48] = 1'b0;
	assign img[19][49] = 1'b0;
	assign img[19][50] = 1'b0;
	assign img[19][51] = 1'b0;
	assign img[19][52] = 1'b0;
	assign img[19][53] = 1'b0;
	assign img[19][54] = 1'b0;
	assign img[19][55] = 1'b0;
	assign img[19][56] = 1'b0;
	assign img[19][57] = 1'b0;
	assign img[19][58] = 1'b0;
	assign img[19][59] = 1'b0;
	assign img[19][60] = 1'b0;
	assign img[19][61] = 1'b0;
	assign img[19][62] = 1'b0;
	assign img[19][63] = 1'b0;
	assign img[20][0] = 1'b0;
	assign img[20][1] = 1'b0;
	assign img[20][2] = 1'b0;
	assign img[20][3] = 1'b0;
	assign img[20][4] = 1'b0;
	assign img[20][5] = 1'b0;
	assign img[20][6] = 1'b0;
	assign img[20][7] = 1'b0;
	assign img[20][8] = 1'b0;
	assign img[20][9] = 1'b0;
	assign img[20][10] = 1'b0;
	assign img[20][11] = 1'b0;
	assign img[20][12] = 1'b0;
	assign img[20][13] = 1'b0;
	assign img[20][14] = 1'b0;
	assign img[20][15] = 1'b0;
	assign img[20][16] = 1'b0;
	assign img[20][17] = 1'b0;
	assign img[20][18] = 1'b0;
	assign img[20][19] = 1'b0;
	assign img[20][20] = 1'b0;
	assign img[20][21] = 1'b0;
	assign img[20][22] = 1'b0;
	assign img[20][23] = 1'b0;
	assign img[20][24] = 1'b0;
	assign img[20][25] = 1'b0;
	assign img[20][26] = 1'b0;
	assign img[20][27] = 1'b0;
	assign img[20][28] = 1'b0;
	assign img[20][29] = 1'b0;
	assign img[20][30] = 1'b0;
	assign img[20][31] = 1'b0;
	assign img[20][32] = 1'b0;
	assign img[20][33] = 1'b0;
	assign img[20][34] = 1'b0;
	assign img[20][35] = 1'b0;
	assign img[20][36] = 1'b0;
	assign img[20][37] = 1'b0;
	assign img[20][38] = 1'b0;
	assign img[20][39] = 1'b0;
	assign img[20][40] = 1'b0;
	assign img[20][41] = 1'b0;
	assign img[20][42] = 1'b0;
	assign img[20][43] = 1'b0;
	assign img[20][44] = 1'b0;
	assign img[20][45] = 1'b0;
	assign img[20][46] = 1'b0;
	assign img[20][47] = 1'b0;
	assign img[20][48] = 1'b0;
	assign img[20][49] = 1'b0;
	assign img[20][50] = 1'b0;
	assign img[20][51] = 1'b0;
	assign img[20][52] = 1'b0;
	assign img[20][53] = 1'b0;
	assign img[20][54] = 1'b0;
	assign img[20][55] = 1'b0;
	assign img[20][56] = 1'b0;
	assign img[20][57] = 1'b0;
	assign img[20][58] = 1'b0;
	assign img[20][59] = 1'b0;
	assign img[20][60] = 1'b0;
	assign img[20][61] = 1'b0;
	assign img[20][62] = 1'b0;
	assign img[20][63] = 1'b0;
	assign img[21][0] = 1'b0;
	assign img[21][1] = 1'b0;
	assign img[21][2] = 1'b0;
	assign img[21][3] = 1'b0;
	assign img[21][4] = 1'b0;
	assign img[21][5] = 1'b0;
	assign img[21][6] = 1'b0;
	assign img[21][7] = 1'b0;
	assign img[21][8] = 1'b0;
	assign img[21][9] = 1'b1;
	assign img[21][10] = 1'b0;
	assign img[21][11] = 1'b0;
	assign img[21][12] = 1'b0;
	assign img[21][13] = 1'b0;
	assign img[21][14] = 1'b0;
	assign img[21][15] = 1'b0;
	assign img[21][16] = 1'b0;
	assign img[21][17] = 1'b0;
	assign img[21][18] = 1'b0;
	assign img[21][19] = 1'b0;
	assign img[21][20] = 1'b0;
	assign img[21][21] = 1'b0;
	assign img[21][22] = 1'b0;
	assign img[21][23] = 1'b0;
	assign img[21][24] = 1'b0;
	assign img[21][25] = 1'b0;
	assign img[21][26] = 1'b0;
	assign img[21][27] = 1'b0;
	assign img[21][28] = 1'b0;
	assign img[21][29] = 1'b0;
	assign img[21][30] = 1'b0;
	assign img[21][31] = 1'b0;
	assign img[21][32] = 1'b0;
	assign img[21][33] = 1'b0;
	assign img[21][34] = 1'b0;
	assign img[21][35] = 1'b0;
	assign img[21][36] = 1'b0;
	assign img[21][37] = 1'b0;
	assign img[21][38] = 1'b0;
	assign img[21][39] = 1'b0;
	assign img[21][40] = 1'b0;
	assign img[21][41] = 1'b0;
	assign img[21][42] = 1'b0;
	assign img[21][43] = 1'b0;
	assign img[21][44] = 1'b0;
	assign img[21][45] = 1'b0;
	assign img[21][46] = 1'b0;
	assign img[21][47] = 1'b0;
	assign img[21][48] = 1'b0;
	assign img[21][49] = 1'b0;
	assign img[21][50] = 1'b0;
	assign img[21][51] = 1'b0;
	assign img[21][52] = 1'b0;
	assign img[21][53] = 1'b0;
	assign img[21][54] = 1'b0;
	assign img[21][55] = 1'b0;
	assign img[21][56] = 1'b0;
	assign img[21][57] = 1'b0;
	assign img[21][58] = 1'b0;
	assign img[21][59] = 1'b0;
	assign img[21][60] = 1'b0;
	assign img[21][61] = 1'b0;
	assign img[21][62] = 1'b0;
	assign img[21][63] = 1'b0;
	assign img[22][0] = 1'b0;
	assign img[22][1] = 1'b0;
	assign img[22][2] = 1'b0;
	assign img[22][3] = 1'b0;
	assign img[22][4] = 1'b0;
	assign img[22][5] = 1'b0;
	assign img[22][6] = 1'b0;
	assign img[22][7] = 1'b0;
	assign img[22][8] = 1'b0;
	assign img[22][9] = 1'b0;
	assign img[22][10] = 1'b0;
	assign img[22][11] = 1'b0;
	assign img[22][12] = 1'b0;
	assign img[22][13] = 1'b0;
	assign img[22][14] = 1'b0;
	assign img[22][15] = 1'b0;
	assign img[22][16] = 1'b0;
	assign img[22][17] = 1'b0;
	assign img[22][18] = 1'b0;
	assign img[22][19] = 1'b0;
	assign img[22][20] = 1'b0;
	assign img[22][21] = 1'b0;
	assign img[22][22] = 1'b0;
	assign img[22][23] = 1'b0;
	assign img[22][24] = 1'b0;
	assign img[22][25] = 1'b0;
	assign img[22][26] = 1'b0;
	assign img[22][27] = 1'b0;
	assign img[22][28] = 1'b0;
	assign img[22][29] = 1'b0;
	assign img[22][30] = 1'b0;
	assign img[22][31] = 1'b0;
	assign img[22][32] = 1'b0;
	assign img[22][33] = 1'b0;
	assign img[22][34] = 1'b0;
	assign img[22][35] = 1'b0;
	assign img[22][36] = 1'b0;
	assign img[22][37] = 1'b0;
	assign img[22][38] = 1'b0;
	assign img[22][39] = 1'b0;
	assign img[22][40] = 1'b0;
	assign img[22][41] = 1'b0;
	assign img[22][42] = 1'b0;
	assign img[22][43] = 1'b0;
	assign img[22][44] = 1'b0;
	assign img[22][45] = 1'b0;
	assign img[22][46] = 1'b0;
	assign img[22][47] = 1'b0;
	assign img[22][48] = 1'b0;
	assign img[22][49] = 1'b0;
	assign img[22][50] = 1'b0;
	assign img[22][51] = 1'b0;
	assign img[22][52] = 1'b0;
	assign img[22][53] = 1'b0;
	assign img[22][54] = 1'b0;
	assign img[22][55] = 1'b0;
	assign img[22][56] = 1'b0;
	assign img[22][57] = 1'b0;
	assign img[22][58] = 1'b0;
	assign img[22][59] = 1'b0;
	assign img[22][60] = 1'b0;
	assign img[22][61] = 1'b0;
	assign img[22][62] = 1'b0;
	assign img[22][63] = 1'b0;
	assign img[23][0] = 1'b0;
	assign img[23][1] = 1'b0;
	assign img[23][2] = 1'b0;
	assign img[23][3] = 1'b0;
	assign img[23][4] = 1'b0;
	assign img[23][5] = 1'b0;
	assign img[23][6] = 1'b0;
	assign img[23][7] = 1'b0;
	assign img[23][8] = 1'b0;
	assign img[23][9] = 1'b0;
	assign img[23][10] = 1'b0;
	assign img[23][11] = 1'b0;
	assign img[23][12] = 1'b0;
	assign img[23][13] = 1'b0;
	assign img[23][14] = 1'b0;
	assign img[23][15] = 1'b0;
	assign img[23][16] = 1'b0;
	assign img[23][17] = 1'b0;
	assign img[23][18] = 1'b0;
	assign img[23][19] = 1'b0;
	assign img[23][20] = 1'b0;
	assign img[23][21] = 1'b0;
	assign img[23][22] = 1'b0;
	assign img[23][23] = 1'b0;
	assign img[23][24] = 1'b0;
	assign img[23][25] = 1'b0;
	assign img[23][26] = 1'b0;
	assign img[23][27] = 1'b0;
	assign img[23][28] = 1'b0;
	assign img[23][29] = 1'b0;
	assign img[23][30] = 1'b0;
	assign img[23][31] = 1'b0;
	assign img[23][32] = 1'b0;
	assign img[23][33] = 1'b0;
	assign img[23][34] = 1'b0;
	assign img[23][35] = 1'b0;
	assign img[23][36] = 1'b0;
	assign img[23][37] = 1'b0;
	assign img[23][38] = 1'b1;
	assign img[23][39] = 1'b0;
	assign img[23][40] = 1'b0;
	assign img[23][41] = 1'b0;
	assign img[23][42] = 1'b0;
	assign img[23][43] = 1'b0;
	assign img[23][44] = 1'b0;
	assign img[23][45] = 1'b0;
	assign img[23][46] = 1'b0;
	assign img[23][47] = 1'b0;
	assign img[23][48] = 1'b0;
	assign img[23][49] = 1'b0;
	assign img[23][50] = 1'b0;
	assign img[23][51] = 1'b0;
	assign img[23][52] = 1'b0;
	assign img[23][53] = 1'b0;
	assign img[23][54] = 1'b0;
	assign img[23][55] = 1'b0;
	assign img[23][56] = 1'b0;
	assign img[23][57] = 1'b0;
	assign img[23][58] = 1'b0;
	assign img[23][59] = 1'b0;
	assign img[23][60] = 1'b0;
	assign img[23][61] = 1'b0;
	assign img[23][62] = 1'b0;
	assign img[23][63] = 1'b0;
	assign img[24][0] = 1'b0;
	assign img[24][1] = 1'b0;
	assign img[24][2] = 1'b0;
	assign img[24][3] = 1'b0;
	assign img[24][4] = 1'b0;
	assign img[24][5] = 1'b0;
	assign img[24][6] = 1'b0;
	assign img[24][7] = 1'b0;
	assign img[24][8] = 1'b0;
	assign img[24][9] = 1'b0;
	assign img[24][10] = 1'b0;
	assign img[24][11] = 1'b0;
	assign img[24][12] = 1'b0;
	assign img[24][13] = 1'b0;
	assign img[24][14] = 1'b0;
	assign img[24][15] = 1'b0;
	assign img[24][16] = 1'b0;
	assign img[24][17] = 1'b0;
	assign img[24][18] = 1'b0;
	assign img[24][19] = 1'b0;
	assign img[24][20] = 1'b0;
	assign img[24][21] = 1'b0;
	assign img[24][22] = 1'b0;
	assign img[24][23] = 1'b0;
	assign img[24][24] = 1'b0;
	assign img[24][25] = 1'b0;
	assign img[24][26] = 1'b0;
	assign img[24][27] = 1'b0;
	assign img[24][28] = 1'b0;
	assign img[24][29] = 1'b0;
	assign img[24][30] = 1'b0;
	assign img[24][31] = 1'b0;
	assign img[24][32] = 1'b0;
	assign img[24][33] = 1'b0;
	assign img[24][34] = 1'b0;
	assign img[24][35] = 1'b0;
	assign img[24][36] = 1'b0;
	assign img[24][37] = 1'b0;
	assign img[24][38] = 1'b0;
	assign img[24][39] = 1'b0;
	assign img[24][40] = 1'b0;
	assign img[24][41] = 1'b0;
	assign img[24][42] = 1'b0;
	assign img[24][43] = 1'b0;
	assign img[24][44] = 1'b0;
	assign img[24][45] = 1'b0;
	assign img[24][46] = 1'b0;
	assign img[24][47] = 1'b0;
	assign img[24][48] = 1'b0;
	assign img[24][49] = 1'b0;
	assign img[24][50] = 1'b0;
	assign img[24][51] = 1'b0;
	assign img[24][52] = 1'b0;
	assign img[24][53] = 1'b0;
	assign img[24][54] = 1'b0;
	assign img[24][55] = 1'b0;
	assign img[24][56] = 1'b0;
	assign img[24][57] = 1'b0;
	assign img[24][58] = 1'b0;
	assign img[24][59] = 1'b0;
	assign img[24][60] = 1'b0;
	assign img[24][61] = 1'b0;
	assign img[24][62] = 1'b0;
	assign img[24][63] = 1'b0;
	assign img[25][0] = 1'b0;
	assign img[25][1] = 1'b0;
	assign img[25][2] = 1'b0;
	assign img[25][3] = 1'b0;
	assign img[25][4] = 1'b0;
	assign img[25][5] = 1'b0;
	assign img[25][6] = 1'b0;
	assign img[25][7] = 1'b0;
	assign img[25][8] = 1'b0;
	assign img[25][9] = 1'b0;
	assign img[25][10] = 1'b0;
	assign img[25][11] = 1'b0;
	assign img[25][12] = 1'b0;
	assign img[25][13] = 1'b0;
	assign img[25][14] = 1'b0;
	assign img[25][15] = 1'b0;
	assign img[25][16] = 1'b0;
	assign img[25][17] = 1'b0;
	assign img[25][18] = 1'b0;
	assign img[25][19] = 1'b0;
	assign img[25][20] = 1'b0;
	assign img[25][21] = 1'b0;
	assign img[25][22] = 1'b0;
	assign img[25][23] = 1'b0;
	assign img[25][24] = 1'b0;
	assign img[25][25] = 1'b0;
	assign img[25][26] = 1'b0;
	assign img[25][27] = 1'b0;
	assign img[25][28] = 1'b0;
	assign img[25][29] = 1'b0;
	assign img[25][30] = 1'b0;
	assign img[25][31] = 1'b0;
	assign img[25][32] = 1'b0;
	assign img[25][33] = 1'b0;
	assign img[25][34] = 1'b0;
	assign img[25][35] = 1'b0;
	assign img[25][36] = 1'b0;
	assign img[25][37] = 1'b0;
	assign img[25][38] = 1'b0;
	assign img[25][39] = 1'b0;
	assign img[25][40] = 1'b0;
	assign img[25][41] = 1'b0;
	assign img[25][42] = 1'b0;
	assign img[25][43] = 1'b0;
	assign img[25][44] = 1'b0;
	assign img[25][45] = 1'b0;
	assign img[25][46] = 1'b0;
	assign img[25][47] = 1'b0;
	assign img[25][48] = 1'b0;
	assign img[25][49] = 1'b0;
	assign img[25][50] = 1'b0;
	assign img[25][51] = 1'b0;
	assign img[25][52] = 1'b0;
	assign img[25][53] = 1'b0;
	assign img[25][54] = 1'b0;
	assign img[25][55] = 1'b0;
	assign img[25][56] = 1'b0;
	assign img[25][57] = 1'b0;
	assign img[25][58] = 1'b0;
	assign img[25][59] = 1'b0;
	assign img[25][60] = 1'b0;
	assign img[25][61] = 1'b0;
	assign img[25][62] = 1'b0;
	assign img[25][63] = 1'b0;
	assign img[26][0] = 1'b0;
	assign img[26][1] = 1'b0;
	assign img[26][2] = 1'b0;
	assign img[26][3] = 1'b0;
	assign img[26][4] = 1'b0;
	assign img[26][5] = 1'b0;
	assign img[26][6] = 1'b0;
	assign img[26][7] = 1'b0;
	assign img[26][8] = 1'b0;
	assign img[26][9] = 1'b0;
	assign img[26][10] = 1'b0;
	assign img[26][11] = 1'b0;
	assign img[26][12] = 1'b0;
	assign img[26][13] = 1'b0;
	assign img[26][14] = 1'b0;
	assign img[26][15] = 1'b0;
	assign img[26][16] = 1'b0;
	assign img[26][17] = 1'b0;
	assign img[26][18] = 1'b0;
	assign img[26][19] = 1'b0;
	assign img[26][20] = 1'b0;
	assign img[26][21] = 1'b0;
	assign img[26][22] = 1'b0;
	assign img[26][23] = 1'b0;
	assign img[26][24] = 1'b0;
	assign img[26][25] = 1'b0;
	assign img[26][26] = 1'b0;
	assign img[26][27] = 1'b0;
	assign img[26][28] = 1'b0;
	assign img[26][29] = 1'b0;
	assign img[26][30] = 1'b0;
	assign img[26][31] = 1'b0;
	assign img[26][32] = 1'b0;
	assign img[26][33] = 1'b0;
	assign img[26][34] = 1'b0;
	assign img[26][35] = 1'b0;
	assign img[26][36] = 1'b0;
	assign img[26][37] = 1'b0;
	assign img[26][38] = 1'b0;
	assign img[26][39] = 1'b0;
	assign img[26][40] = 1'b0;
	assign img[26][41] = 1'b0;
	assign img[26][42] = 1'b0;
	assign img[26][43] = 1'b0;
	assign img[26][44] = 1'b0;
	assign img[26][45] = 1'b0;
	assign img[26][46] = 1'b0;
	assign img[26][47] = 1'b0;
	assign img[26][48] = 1'b0;
	assign img[26][49] = 1'b0;
	assign img[26][50] = 1'b0;
	assign img[26][51] = 1'b0;
	assign img[26][52] = 1'b0;
	assign img[26][53] = 1'b0;
	assign img[26][54] = 1'b0;
	assign img[26][55] = 1'b0;
	assign img[26][56] = 1'b0;
	assign img[26][57] = 1'b0;
	assign img[26][58] = 1'b0;
	assign img[26][59] = 1'b0;
	assign img[26][60] = 1'b0;
	assign img[26][61] = 1'b0;
	assign img[26][62] = 1'b0;
	assign img[26][63] = 1'b0;
	assign img[27][0] = 1'b0;
	assign img[27][1] = 1'b0;
	assign img[27][2] = 1'b0;
	assign img[27][3] = 1'b0;
	assign img[27][4] = 1'b0;
	assign img[27][5] = 1'b0;
	assign img[27][6] = 1'b0;
	assign img[27][7] = 1'b0;
	assign img[27][8] = 1'b0;
	assign img[27][9] = 1'b0;
	assign img[27][10] = 1'b0;
	assign img[27][11] = 1'b0;
	assign img[27][12] = 1'b0;
	assign img[27][13] = 1'b0;
	assign img[27][14] = 1'b0;
	assign img[27][15] = 1'b0;
	assign img[27][16] = 1'b0;
	assign img[27][17] = 1'b0;
	assign img[27][18] = 1'b0;
	assign img[27][19] = 1'b0;
	assign img[27][20] = 1'b0;
	assign img[27][21] = 1'b0;
	assign img[27][22] = 1'b0;
	assign img[27][23] = 1'b0;
	assign img[27][24] = 1'b0;
	assign img[27][25] = 1'b0;
	assign img[27][26] = 1'b0;
	assign img[27][27] = 1'b0;
	assign img[27][28] = 1'b0;
	assign img[27][29] = 1'b0;
	assign img[27][30] = 1'b0;
	assign img[27][31] = 1'b0;
	assign img[27][32] = 1'b0;
	assign img[27][33] = 1'b0;
	assign img[27][34] = 1'b0;
	assign img[27][35] = 1'b0;
	assign img[27][36] = 1'b0;
	assign img[27][37] = 1'b0;
	assign img[27][38] = 1'b0;
	assign img[27][39] = 1'b0;
	assign img[27][40] = 1'b0;
	assign img[27][41] = 1'b0;
	assign img[27][42] = 1'b0;
	assign img[27][43] = 1'b0;
	assign img[27][44] = 1'b0;
	assign img[27][45] = 1'b0;
	assign img[27][46] = 1'b0;
	assign img[27][47] = 1'b0;
	assign img[27][48] = 1'b0;
	assign img[27][49] = 1'b0;
	assign img[27][50] = 1'b0;
	assign img[27][51] = 1'b0;
	assign img[27][52] = 1'b0;
	assign img[27][53] = 1'b0;
	assign img[27][54] = 1'b0;
	assign img[27][55] = 1'b0;
	assign img[27][56] = 1'b0;
	assign img[27][57] = 1'b0;
	assign img[27][58] = 1'b0;
	assign img[27][59] = 1'b0;
	assign img[27][60] = 1'b0;
	assign img[27][61] = 1'b0;
	assign img[27][62] = 1'b0;
	assign img[27][63] = 1'b0;
	assign img[28][0] = 1'b0;
	assign img[28][1] = 1'b0;
	assign img[28][2] = 1'b0;
	assign img[28][3] = 1'b0;
	assign img[28][4] = 1'b0;
	assign img[28][5] = 1'b0;
	assign img[28][6] = 1'b0;
	assign img[28][7] = 1'b0;
	assign img[28][8] = 1'b0;
	assign img[28][9] = 1'b0;
	assign img[28][10] = 1'b0;
	assign img[28][11] = 1'b0;
	assign img[28][12] = 1'b0;
	assign img[28][13] = 1'b0;
	assign img[28][14] = 1'b0;
	assign img[28][15] = 1'b0;
	assign img[28][16] = 1'b0;
	assign img[28][17] = 1'b0;
	assign img[28][18] = 1'b0;
	assign img[28][19] = 1'b0;
	assign img[28][20] = 1'b0;
	assign img[28][21] = 1'b0;
	assign img[28][22] = 1'b0;
	assign img[28][23] = 1'b0;
	assign img[28][24] = 1'b0;
	assign img[28][25] = 1'b0;
	assign img[28][26] = 1'b0;
	assign img[28][27] = 1'b0;
	assign img[28][28] = 1'b0;
	assign img[28][29] = 1'b0;
	assign img[28][30] = 1'b0;
	assign img[28][31] = 1'b0;
	assign img[28][32] = 1'b0;
	assign img[28][33] = 1'b0;
	assign img[28][34] = 1'b0;
	assign img[28][35] = 1'b0;
	assign img[28][36] = 1'b0;
	assign img[28][37] = 1'b0;
	assign img[28][38] = 1'b0;
	assign img[28][39] = 1'b0;
	assign img[28][40] = 1'b0;
	assign img[28][41] = 1'b0;
	assign img[28][42] = 1'b0;
	assign img[28][43] = 1'b0;
	assign img[28][44] = 1'b0;
	assign img[28][45] = 1'b0;
	assign img[28][46] = 1'b0;
	assign img[28][47] = 1'b0;
	assign img[28][48] = 1'b0;
	assign img[28][49] = 1'b0;
	assign img[28][50] = 1'b0;
	assign img[28][51] = 1'b0;
	assign img[28][52] = 1'b0;
	assign img[28][53] = 1'b0;
	assign img[28][54] = 1'b0;
	assign img[28][55] = 1'b0;
	assign img[28][56] = 1'b0;
	assign img[28][57] = 1'b0;
	assign img[28][58] = 1'b0;
	assign img[28][59] = 1'b1;
	assign img[28][60] = 1'b0;
	assign img[28][61] = 1'b0;
	assign img[28][62] = 1'b0;
	assign img[28][63] = 1'b0;
	assign img[29][0] = 1'b0;
	assign img[29][1] = 1'b0;
	assign img[29][2] = 1'b0;
	assign img[29][3] = 1'b0;
	assign img[29][4] = 1'b0;
	assign img[29][5] = 1'b0;
	assign img[29][6] = 1'b0;
	assign img[29][7] = 1'b0;
	assign img[29][8] = 1'b0;
	assign img[29][9] = 1'b0;
	assign img[29][10] = 1'b0;
	assign img[29][11] = 1'b0;
	assign img[29][12] = 1'b0;
	assign img[29][13] = 1'b0;
	assign img[29][14] = 1'b0;
	assign img[29][15] = 1'b0;
	assign img[29][16] = 1'b0;
	assign img[29][17] = 1'b0;
	assign img[29][18] = 1'b0;
	assign img[29][19] = 1'b0;
	assign img[29][20] = 1'b0;
	assign img[29][21] = 1'b0;
	assign img[29][22] = 1'b0;
	assign img[29][23] = 1'b0;
	assign img[29][24] = 1'b0;
	assign img[29][25] = 1'b0;
	assign img[29][26] = 1'b0;
	assign img[29][27] = 1'b0;
	assign img[29][28] = 1'b0;
	assign img[29][29] = 1'b0;
	assign img[29][30] = 1'b0;
	assign img[29][31] = 1'b0;
	assign img[29][32] = 1'b0;
	assign img[29][33] = 1'b1;
	assign img[29][34] = 1'b0;
	assign img[29][35] = 1'b0;
	assign img[29][36] = 1'b0;
	assign img[29][37] = 1'b0;
	assign img[29][38] = 1'b0;
	assign img[29][39] = 1'b0;
	assign img[29][40] = 1'b0;
	assign img[29][41] = 1'b0;
	assign img[29][42] = 1'b0;
	assign img[29][43] = 1'b0;
	assign img[29][44] = 1'b0;
	assign img[29][45] = 1'b0;
	assign img[29][46] = 1'b0;
	assign img[29][47] = 1'b0;
	assign img[29][48] = 1'b0;
	assign img[29][49] = 1'b0;
	assign img[29][50] = 1'b1;
	assign img[29][51] = 1'b0;
	assign img[29][52] = 1'b0;
	assign img[29][53] = 1'b0;
	assign img[29][54] = 1'b0;
	assign img[29][55] = 1'b1;
	assign img[29][56] = 1'b0;
	assign img[29][57] = 1'b0;
	assign img[29][58] = 1'b0;
	assign img[29][59] = 1'b0;
	assign img[29][60] = 1'b0;
	assign img[29][61] = 1'b0;
	assign img[29][62] = 1'b0;
	assign img[29][63] = 1'b0;
	assign img[30][0] = 1'b0;
	assign img[30][1] = 1'b0;
	assign img[30][2] = 1'b0;
	assign img[30][3] = 1'b0;
	assign img[30][4] = 1'b0;
	assign img[30][5] = 1'b0;
	assign img[30][6] = 1'b0;
	assign img[30][7] = 1'b0;
	assign img[30][8] = 1'b0;
	assign img[30][9] = 1'b0;
	assign img[30][10] = 1'b1;
	assign img[30][11] = 1'b0;
	assign img[30][12] = 1'b0;
	assign img[30][13] = 1'b0;
	assign img[30][14] = 1'b1;
	assign img[30][15] = 1'b0;
	assign img[30][16] = 1'b0;
	assign img[30][17] = 1'b0;
	assign img[30][18] = 1'b0;
	assign img[30][19] = 1'b0;
	assign img[30][20] = 1'b0;
	assign img[30][21] = 1'b0;
	assign img[30][22] = 1'b0;
	assign img[30][23] = 1'b0;
	assign img[30][24] = 1'b0;
	assign img[30][25] = 1'b0;
	assign img[30][26] = 1'b0;
	assign img[30][27] = 1'b0;
	assign img[30][28] = 1'b0;
	assign img[30][29] = 1'b0;
	assign img[30][30] = 1'b0;
	assign img[30][31] = 1'b0;
	assign img[30][32] = 1'b0;
	assign img[30][33] = 1'b0;
	assign img[30][34] = 1'b0;
	assign img[30][35] = 1'b1;
	assign img[30][36] = 1'b0;
	assign img[30][37] = 1'b0;
	assign img[30][38] = 1'b0;
	assign img[30][39] = 1'b0;
	assign img[30][40] = 1'b0;
	assign img[30][41] = 1'b0;
	assign img[30][42] = 1'b0;
	assign img[30][43] = 1'b0;
	assign img[30][44] = 1'b0;
	assign img[30][45] = 1'b0;
	assign img[30][46] = 1'b0;
	assign img[30][47] = 1'b0;
	assign img[30][48] = 1'b0;
	assign img[30][49] = 1'b0;
	assign img[30][50] = 1'b0;
	assign img[30][51] = 1'b0;
	assign img[30][52] = 1'b0;
	assign img[30][53] = 1'b0;
	assign img[30][54] = 1'b0;
	assign img[30][55] = 1'b0;
	assign img[30][56] = 1'b0;
	assign img[30][57] = 1'b0;
	assign img[30][58] = 1'b0;
	assign img[30][59] = 1'b0;
	assign img[30][60] = 1'b0;
	assign img[30][61] = 1'b0;
	assign img[30][62] = 1'b0;
	assign img[30][63] = 1'b0;
	assign img[31][0] = 1'b0;
	assign img[31][1] = 1'b0;
	assign img[31][2] = 1'b0;
	assign img[31][3] = 1'b0;
	assign img[31][4] = 1'b0;
	assign img[31][5] = 1'b0;
	assign img[31][6] = 1'b0;
	assign img[31][7] = 1'b0;
	assign img[31][8] = 1'b0;
	assign img[31][9] = 1'b0;
	assign img[31][10] = 1'b0;
	assign img[31][11] = 1'b0;
	assign img[31][12] = 1'b0;
	assign img[31][13] = 1'b0;
	assign img[31][14] = 1'b0;
	assign img[31][15] = 1'b0;
	assign img[31][16] = 1'b0;
	assign img[31][17] = 1'b0;
	assign img[31][18] = 1'b0;
	assign img[31][19] = 1'b0;
	assign img[31][20] = 1'b0;
	assign img[31][21] = 1'b0;
	assign img[31][22] = 1'b0;
	assign img[31][23] = 1'b0;
	assign img[31][24] = 1'b0;
	assign img[31][25] = 1'b0;
	assign img[31][26] = 1'b0;
	assign img[31][27] = 1'b1;
	assign img[31][28] = 1'b0;
	assign img[31][29] = 1'b0;
	assign img[31][30] = 1'b0;
	assign img[31][31] = 1'b0;
	assign img[31][32] = 1'b0;
	assign img[31][33] = 1'b0;
	assign img[31][34] = 1'b0;
	assign img[31][35] = 1'b0;
	assign img[31][36] = 1'b0;
	assign img[31][37] = 1'b0;
	assign img[31][38] = 1'b0;
	assign img[31][39] = 1'b0;
	assign img[31][40] = 1'b0;
	assign img[31][41] = 1'b0;
	assign img[31][42] = 1'b0;
	assign img[31][43] = 1'b0;
	assign img[31][44] = 1'b0;
	assign img[31][45] = 1'b0;
	assign img[31][46] = 1'b0;
	assign img[31][47] = 1'b0;
	assign img[31][48] = 1'b0;
	assign img[31][49] = 1'b0;
	assign img[31][50] = 1'b0;
	assign img[31][51] = 1'b0;
	assign img[31][52] = 1'b0;
	assign img[31][53] = 1'b0;
	assign img[31][54] = 1'b0;
	assign img[31][55] = 1'b0;
	assign img[31][56] = 1'b0;
	assign img[31][57] = 1'b0;
	assign img[31][58] = 1'b0;
	assign img[31][59] = 1'b0;
	assign img[31][60] = 1'b0;
	assign img[31][61] = 1'b0;
	assign img[31][62] = 1'b0;
	assign img[31][63] = 1'b0;
	assign img[32][0] = 1'b0;
	assign img[32][1] = 1'b0;
	assign img[32][2] = 1'b0;
	assign img[32][3] = 1'b0;
	assign img[32][4] = 1'b0;
	assign img[32][5] = 1'b0;
	assign img[32][6] = 1'b0;
	assign img[32][7] = 1'b0;
	assign img[32][8] = 1'b0;
	assign img[32][9] = 1'b0;
	assign img[32][10] = 1'b0;
	assign img[32][11] = 1'b0;
	assign img[32][12] = 1'b0;
	assign img[32][13] = 1'b0;
	assign img[32][14] = 1'b0;
	assign img[32][15] = 1'b0;
	assign img[32][16] = 1'b0;
	assign img[32][17] = 1'b0;
	assign img[32][18] = 1'b0;
	assign img[32][19] = 1'b1;
	assign img[32][20] = 1'b0;
	assign img[32][21] = 1'b0;
	assign img[32][22] = 1'b0;
	assign img[32][23] = 1'b0;
	assign img[32][24] = 1'b0;
	assign img[32][25] = 1'b0;
	assign img[32][26] = 1'b0;
	assign img[32][27] = 1'b0;
	assign img[32][28] = 1'b0;
	assign img[32][29] = 1'b0;
	assign img[32][30] = 1'b0;
	assign img[32][31] = 1'b0;
	assign img[32][32] = 1'b0;
	assign img[32][33] = 1'b0;
	assign img[32][34] = 1'b0;
	assign img[32][35] = 1'b0;
	assign img[32][36] = 1'b0;
	assign img[32][37] = 1'b0;
	assign img[32][38] = 1'b0;
	assign img[32][39] = 1'b0;
	assign img[32][40] = 1'b0;
	assign img[32][41] = 1'b0;
	assign img[32][42] = 1'b0;
	assign img[32][43] = 1'b0;
	assign img[32][44] = 1'b0;
	assign img[32][45] = 1'b0;
	assign img[32][46] = 1'b0;
	assign img[32][47] = 1'b0;
	assign img[32][48] = 1'b0;
	assign img[32][49] = 1'b0;
	assign img[32][50] = 1'b0;
	assign img[32][51] = 1'b0;
	assign img[32][52] = 1'b0;
	assign img[32][53] = 1'b0;
	assign img[32][54] = 1'b0;
	assign img[32][55] = 1'b0;
	assign img[32][56] = 1'b0;
	assign img[32][57] = 1'b0;
	assign img[32][58] = 1'b0;
	assign img[32][59] = 1'b0;
	assign img[32][60] = 1'b0;
	assign img[32][61] = 1'b0;
	assign img[32][62] = 1'b0;
	assign img[32][63] = 1'b0;
	assign img[33][0] = 1'b0;
	assign img[33][1] = 1'b0;
	assign img[33][2] = 1'b0;
	assign img[33][3] = 1'b0;
	assign img[33][4] = 1'b0;
	assign img[33][5] = 1'b0;
	assign img[33][6] = 1'b0;
	assign img[33][7] = 1'b0;
	assign img[33][8] = 1'b0;
	assign img[33][9] = 1'b0;
	assign img[33][10] = 1'b0;
	assign img[33][11] = 1'b0;
	assign img[33][12] = 1'b0;
	assign img[33][13] = 1'b0;
	assign img[33][14] = 1'b0;
	assign img[33][15] = 1'b0;
	assign img[33][16] = 1'b0;
	assign img[33][17] = 1'b0;
	assign img[33][18] = 1'b0;
	assign img[33][19] = 1'b0;
	assign img[33][20] = 1'b0;
	assign img[33][21] = 1'b0;
	assign img[33][22] = 1'b0;
	assign img[33][23] = 1'b0;
	assign img[33][24] = 1'b0;
	assign img[33][25] = 1'b0;
	assign img[33][26] = 1'b0;
	assign img[33][27] = 1'b1;
	assign img[33][28] = 1'b0;
	assign img[33][29] = 1'b0;
	assign img[33][30] = 1'b0;
	assign img[33][31] = 1'b0;
	assign img[33][32] = 1'b0;
	assign img[33][33] = 1'b0;
	assign img[33][34] = 1'b0;
	assign img[33][35] = 1'b0;
	assign img[33][36] = 1'b0;
	assign img[33][37] = 1'b0;
	assign img[33][38] = 1'b0;
	assign img[33][39] = 1'b1;
	assign img[33][40] = 1'b0;
	assign img[33][41] = 1'b0;
	assign img[33][42] = 1'b0;
	assign img[33][43] = 1'b0;
	assign img[33][44] = 1'b0;
	assign img[33][45] = 1'b0;
	assign img[33][46] = 1'b0;
	assign img[33][47] = 1'b0;
	assign img[33][48] = 1'b0;
	assign img[33][49] = 1'b0;
	assign img[33][50] = 1'b0;
	assign img[33][51] = 1'b0;
	assign img[33][52] = 1'b0;
	assign img[33][53] = 1'b0;
	assign img[33][54] = 1'b0;
	assign img[33][55] = 1'b0;
	assign img[33][56] = 1'b0;
	assign img[33][57] = 1'b0;
	assign img[33][58] = 1'b0;
	assign img[33][59] = 1'b0;
	assign img[33][60] = 1'b1;
	assign img[33][61] = 1'b0;
	assign img[33][62] = 1'b0;
	assign img[33][63] = 1'b0;
	assign img[34][0] = 1'b0;
	assign img[34][1] = 1'b0;
	assign img[34][2] = 1'b0;
	assign img[34][3] = 1'b0;
	assign img[34][4] = 1'b0;
	assign img[34][5] = 1'b0;
	assign img[34][6] = 1'b0;
	assign img[34][7] = 1'b0;
	assign img[34][8] = 1'b0;
	assign img[34][9] = 1'b0;
	assign img[34][10] = 1'b0;
	assign img[34][11] = 1'b0;
	assign img[34][12] = 1'b0;
	assign img[34][13] = 1'b0;
	assign img[34][14] = 1'b0;
	assign img[34][15] = 1'b0;
	assign img[34][16] = 1'b0;
	assign img[34][17] = 1'b0;
	assign img[34][18] = 1'b0;
	assign img[34][19] = 1'b0;
	assign img[34][20] = 1'b0;
	assign img[34][21] = 1'b0;
	assign img[34][22] = 1'b0;
	assign img[34][23] = 1'b0;
	assign img[34][24] = 1'b0;
	assign img[34][25] = 1'b0;
	assign img[34][26] = 1'b0;
	assign img[34][27] = 1'b0;
	assign img[34][28] = 1'b0;
	assign img[34][29] = 1'b0;
	assign img[34][30] = 1'b0;
	assign img[34][31] = 1'b0;
	assign img[34][32] = 1'b0;
	assign img[34][33] = 1'b0;
	assign img[34][34] = 1'b0;
	assign img[34][35] = 1'b0;
	assign img[34][36] = 1'b0;
	assign img[34][37] = 1'b0;
	assign img[34][38] = 1'b0;
	assign img[34][39] = 1'b0;
	assign img[34][40] = 1'b0;
	assign img[34][41] = 1'b0;
	assign img[34][42] = 1'b0;
	assign img[34][43] = 1'b0;
	assign img[34][44] = 1'b0;
	assign img[34][45] = 1'b0;
	assign img[34][46] = 1'b0;
	assign img[34][47] = 1'b0;
	assign img[34][48] = 1'b0;
	assign img[34][49] = 1'b0;
	assign img[34][50] = 1'b0;
	assign img[34][51] = 1'b0;
	assign img[34][52] = 1'b0;
	assign img[34][53] = 1'b0;
	assign img[34][54] = 1'b0;
	assign img[34][55] = 1'b0;
	assign img[34][56] = 1'b1;
	assign img[34][57] = 1'b0;
	assign img[34][58] = 1'b0;
	assign img[34][59] = 1'b0;
	assign img[34][60] = 1'b0;
	assign img[34][61] = 1'b0;
	assign img[34][62] = 1'b0;
	assign img[34][63] = 1'b0;
	assign img[35][0] = 1'b0;
	assign img[35][1] = 1'b0;
	assign img[35][2] = 1'b0;
	assign img[35][3] = 1'b0;
	assign img[35][4] = 1'b0;
	assign img[35][5] = 1'b0;
	assign img[35][6] = 1'b0;
	assign img[35][7] = 1'b0;
	assign img[35][8] = 1'b0;
	assign img[35][9] = 1'b0;
	assign img[35][10] = 1'b0;
	assign img[35][11] = 1'b0;
	assign img[35][12] = 1'b0;
	assign img[35][13] = 1'b1;
	assign img[35][14] = 1'b0;
	assign img[35][15] = 1'b0;
	assign img[35][16] = 1'b0;
	assign img[35][17] = 1'b0;
	assign img[35][18] = 1'b0;
	assign img[35][19] = 1'b0;
	assign img[35][20] = 1'b0;
	assign img[35][21] = 1'b0;
	assign img[35][22] = 1'b0;
	assign img[35][23] = 1'b0;
	assign img[35][24] = 1'b0;
	assign img[35][25] = 1'b0;
	assign img[35][26] = 1'b0;
	assign img[35][27] = 1'b0;
	assign img[35][28] = 1'b0;
	assign img[35][29] = 1'b0;
	assign img[35][30] = 1'b0;
	assign img[35][31] = 1'b0;
	assign img[35][32] = 1'b0;
	assign img[35][33] = 1'b0;
	assign img[35][34] = 1'b0;
	assign img[35][35] = 1'b0;
	assign img[35][36] = 1'b0;
	assign img[35][37] = 1'b0;
	assign img[35][38] = 1'b0;
	assign img[35][39] = 1'b0;
	assign img[35][40] = 1'b0;
	assign img[35][41] = 1'b0;
	assign img[35][42] = 1'b0;
	assign img[35][43] = 1'b0;
	assign img[35][44] = 1'b0;
	assign img[35][45] = 1'b0;
	assign img[35][46] = 1'b0;
	assign img[35][47] = 1'b0;
	assign img[35][48] = 1'b0;
	assign img[35][49] = 1'b0;
	assign img[35][50] = 1'b0;
	assign img[35][51] = 1'b0;
	assign img[35][52] = 1'b0;
	assign img[35][53] = 1'b0;
	assign img[35][54] = 1'b0;
	assign img[35][55] = 1'b0;
	assign img[35][56] = 1'b0;
	assign img[35][57] = 1'b0;
	assign img[35][58] = 1'b0;
	assign img[35][59] = 1'b0;
	assign img[35][60] = 1'b0;
	assign img[35][61] = 1'b0;
	assign img[35][62] = 1'b0;
	assign img[35][63] = 1'b0;
	assign img[36][0] = 1'b0;
	assign img[36][1] = 1'b0;
	assign img[36][2] = 1'b0;
	assign img[36][3] = 1'b0;
	assign img[36][4] = 1'b0;
	assign img[36][5] = 1'b0;
	assign img[36][6] = 1'b1;
	assign img[36][7] = 1'b0;
	assign img[36][8] = 1'b0;
	assign img[36][9] = 1'b0;
	assign img[36][10] = 1'b0;
	assign img[36][11] = 1'b0;
	assign img[36][12] = 1'b0;
	assign img[36][13] = 1'b0;
	assign img[36][14] = 1'b0;
	assign img[36][15] = 1'b0;
	assign img[36][16] = 1'b0;
	assign img[36][17] = 1'b1;
	assign img[36][18] = 1'b0;
	assign img[36][19] = 1'b0;
	assign img[36][20] = 1'b0;
	assign img[36][21] = 1'b0;
	assign img[36][22] = 1'b0;
	assign img[36][23] = 1'b0;
	assign img[36][24] = 1'b0;
	assign img[36][25] = 1'b0;
	assign img[36][26] = 1'b0;
	assign img[36][27] = 1'b0;
	assign img[36][28] = 1'b0;
	assign img[36][29] = 1'b0;
	assign img[36][30] = 1'b0;
	assign img[36][31] = 1'b0;
	assign img[36][32] = 1'b0;
	assign img[36][33] = 1'b0;
	assign img[36][34] = 1'b0;
	assign img[36][35] = 1'b0;
	assign img[36][36] = 1'b0;
	assign img[36][37] = 1'b0;
	assign img[36][38] = 1'b0;
	assign img[36][39] = 1'b0;
	assign img[36][40] = 1'b0;
	assign img[36][41] = 1'b0;
	assign img[36][42] = 1'b0;
	assign img[36][43] = 1'b0;
	assign img[36][44] = 1'b0;
	assign img[36][45] = 1'b0;
	assign img[36][46] = 1'b0;
	assign img[36][47] = 1'b0;
	assign img[36][48] = 1'b0;
	assign img[36][49] = 1'b0;
	assign img[36][50] = 1'b0;
	assign img[36][51] = 1'b0;
	assign img[36][52] = 1'b0;
	assign img[36][53] = 1'b0;
	assign img[36][54] = 1'b0;
	assign img[36][55] = 1'b0;
	assign img[36][56] = 1'b0;
	assign img[36][57] = 1'b0;
	assign img[36][58] = 1'b0;
	assign img[36][59] = 1'b0;
	assign img[36][60] = 1'b0;
	assign img[36][61] = 1'b0;
	assign img[36][62] = 1'b0;
	assign img[36][63] = 1'b0;
	assign img[37][0] = 1'b0;
	assign img[37][1] = 1'b0;
	assign img[37][2] = 1'b0;
	assign img[37][3] = 1'b0;
	assign img[37][4] = 1'b0;
	assign img[37][5] = 1'b0;
	assign img[37][6] = 1'b0;
	assign img[37][7] = 1'b0;
	assign img[37][8] = 1'b0;
	assign img[37][9] = 1'b0;
	assign img[37][10] = 1'b0;
	assign img[37][11] = 1'b0;
	assign img[37][12] = 1'b0;
	assign img[37][13] = 1'b0;
	assign img[37][14] = 1'b0;
	assign img[37][15] = 1'b0;
	assign img[37][16] = 1'b1;
	assign img[37][17] = 1'b0;
	assign img[37][18] = 1'b0;
	assign img[37][19] = 1'b0;
	assign img[37][20] = 1'b0;
	assign img[37][21] = 1'b0;
	assign img[37][22] = 1'b0;
	assign img[37][23] = 1'b0;
	assign img[37][24] = 1'b0;
	assign img[37][25] = 1'b0;
	assign img[37][26] = 1'b0;
	assign img[37][27] = 1'b0;
	assign img[37][28] = 1'b0;
	assign img[37][29] = 1'b0;
	assign img[37][30] = 1'b0;
	assign img[37][31] = 1'b0;
	assign img[37][32] = 1'b0;
	assign img[37][33] = 1'b0;
	assign img[37][34] = 1'b0;
	assign img[37][35] = 1'b0;
	assign img[37][36] = 1'b0;
	assign img[37][37] = 1'b0;
	assign img[37][38] = 1'b0;
	assign img[37][39] = 1'b0;
	assign img[37][40] = 1'b0;
	assign img[37][41] = 1'b0;
	assign img[37][42] = 1'b0;
	assign img[37][43] = 1'b0;
	assign img[37][44] = 1'b0;
	assign img[37][45] = 1'b0;
	assign img[37][46] = 1'b0;
	assign img[37][47] = 1'b0;
	assign img[37][48] = 1'b0;
	assign img[37][49] = 1'b0;
	assign img[37][50] = 1'b0;
	assign img[37][51] = 1'b0;
	assign img[37][52] = 1'b0;
	assign img[37][53] = 1'b0;
	assign img[37][54] = 1'b0;
	assign img[37][55] = 1'b0;
	assign img[37][56] = 1'b0;
	assign img[37][57] = 1'b0;
	assign img[37][58] = 1'b0;
	assign img[37][59] = 1'b0;
	assign img[37][60] = 1'b0;
	assign img[37][61] = 1'b0;
	assign img[37][62] = 1'b0;
	assign img[37][63] = 1'b0;
	assign img[38][0] = 1'b0;
	assign img[38][1] = 1'b0;
	assign img[38][2] = 1'b0;
	assign img[38][3] = 1'b0;
	assign img[38][4] = 1'b0;
	assign img[38][5] = 1'b0;
	assign img[38][6] = 1'b0;
	assign img[38][7] = 1'b0;
	assign img[38][8] = 1'b0;
	assign img[38][9] = 1'b0;
	assign img[38][10] = 1'b0;
	assign img[38][11] = 1'b0;
	assign img[38][12] = 1'b0;
	assign img[38][13] = 1'b0;
	assign img[38][14] = 1'b0;
	assign img[38][15] = 1'b0;
	assign img[38][16] = 1'b0;
	assign img[38][17] = 1'b0;
	assign img[38][18] = 1'b0;
	assign img[38][19] = 1'b0;
	assign img[38][20] = 1'b0;
	assign img[38][21] = 1'b0;
	assign img[38][22] = 1'b0;
	assign img[38][23] = 1'b0;
	assign img[38][24] = 1'b0;
	assign img[38][25] = 1'b0;
	assign img[38][26] = 1'b0;
	assign img[38][27] = 1'b0;
	assign img[38][28] = 1'b0;
	assign img[38][29] = 1'b0;
	assign img[38][30] = 1'b0;
	assign img[38][31] = 1'b0;
	assign img[38][32] = 1'b0;
	assign img[38][33] = 1'b0;
	assign img[38][34] = 1'b0;
	assign img[38][35] = 1'b0;
	assign img[38][36] = 1'b0;
	assign img[38][37] = 1'b0;
	assign img[38][38] = 1'b0;
	assign img[38][39] = 1'b0;
	assign img[38][40] = 1'b0;
	assign img[38][41] = 1'b0;
	assign img[38][42] = 1'b0;
	assign img[38][43] = 1'b0;
	assign img[38][44] = 1'b0;
	assign img[38][45] = 1'b0;
	assign img[38][46] = 1'b0;
	assign img[38][47] = 1'b0;
	assign img[38][48] = 1'b0;
	assign img[38][49] = 1'b0;
	assign img[38][50] = 1'b0;
	assign img[38][51] = 1'b0;
	assign img[38][52] = 1'b0;
	assign img[38][53] = 1'b0;
	assign img[38][54] = 1'b0;
	assign img[38][55] = 1'b0;
	assign img[38][56] = 1'b0;
	assign img[38][57] = 1'b0;
	assign img[38][58] = 1'b0;
	assign img[38][59] = 1'b0;
	assign img[38][60] = 1'b0;
	assign img[38][61] = 1'b0;
	assign img[38][62] = 1'b0;
	assign img[38][63] = 1'b0;
	assign img[39][0] = 1'b0;
	assign img[39][1] = 1'b0;
	assign img[39][2] = 1'b0;
	assign img[39][3] = 1'b0;
	assign img[39][4] = 1'b0;
	assign img[39][5] = 1'b0;
	assign img[39][6] = 1'b0;
	assign img[39][7] = 1'b0;
	assign img[39][8] = 1'b0;
	assign img[39][9] = 1'b0;
	assign img[39][10] = 1'b0;
	assign img[39][11] = 1'b0;
	assign img[39][12] = 1'b0;
	assign img[39][13] = 1'b0;
	assign img[39][14] = 1'b0;
	assign img[39][15] = 1'b0;
	assign img[39][16] = 1'b0;
	assign img[39][17] = 1'b0;
	assign img[39][18] = 1'b0;
	assign img[39][19] = 1'b0;
	assign img[39][20] = 1'b0;
	assign img[39][21] = 1'b0;
	assign img[39][22] = 1'b0;
	assign img[39][23] = 1'b0;
	assign img[39][24] = 1'b0;
	assign img[39][25] = 1'b0;
	assign img[39][26] = 1'b0;
	assign img[39][27] = 1'b0;
	assign img[39][28] = 1'b0;
	assign img[39][29] = 1'b0;
	assign img[39][30] = 1'b0;
	assign img[39][31] = 1'b0;
	assign img[39][32] = 1'b0;
	assign img[39][33] = 1'b0;
	assign img[39][34] = 1'b0;
	assign img[39][35] = 1'b0;
	assign img[39][36] = 1'b0;
	assign img[39][37] = 1'b0;
	assign img[39][38] = 1'b0;
	assign img[39][39] = 1'b0;
	assign img[39][40] = 1'b0;
	assign img[39][41] = 1'b0;
	assign img[39][42] = 1'b0;
	assign img[39][43] = 1'b0;
	assign img[39][44] = 1'b0;
	assign img[39][45] = 1'b0;
	assign img[39][46] = 1'b0;
	assign img[39][47] = 1'b0;
	assign img[39][48] = 1'b0;
	assign img[39][49] = 1'b0;
	assign img[39][50] = 1'b0;
	assign img[39][51] = 1'b0;
	assign img[39][52] = 1'b0;
	assign img[39][53] = 1'b0;
	assign img[39][54] = 1'b0;
	assign img[39][55] = 1'b0;
	assign img[39][56] = 1'b0;
	assign img[39][57] = 1'b0;
	assign img[39][58] = 1'b0;
	assign img[39][59] = 1'b0;
	assign img[39][60] = 1'b0;
	assign img[39][61] = 1'b0;
	assign img[39][62] = 1'b0;
	assign img[39][63] = 1'b0;
	assign img[40][0] = 1'b0;
	assign img[40][1] = 1'b0;
	assign img[40][2] = 1'b0;
	assign img[40][3] = 1'b0;
	assign img[40][4] = 1'b0;
	assign img[40][5] = 1'b0;
	assign img[40][6] = 1'b0;
	assign img[40][7] = 1'b0;
	assign img[40][8] = 1'b0;
	assign img[40][9] = 1'b0;
	assign img[40][10] = 1'b0;
	assign img[40][11] = 1'b0;
	assign img[40][12] = 1'b0;
	assign img[40][13] = 1'b0;
	assign img[40][14] = 1'b0;
	assign img[40][15] = 1'b0;
	assign img[40][16] = 1'b0;
	assign img[40][17] = 1'b0;
	assign img[40][18] = 1'b0;
	assign img[40][19] = 1'b0;
	assign img[40][20] = 1'b0;
	assign img[40][21] = 1'b0;
	assign img[40][22] = 1'b0;
	assign img[40][23] = 1'b0;
	assign img[40][24] = 1'b0;
	assign img[40][25] = 1'b0;
	assign img[40][26] = 1'b0;
	assign img[40][27] = 1'b0;
	assign img[40][28] = 1'b0;
	assign img[40][29] = 1'b0;
	assign img[40][30] = 1'b0;
	assign img[40][31] = 1'b0;
	assign img[40][32] = 1'b0;
	assign img[40][33] = 1'b0;
	assign img[40][34] = 1'b0;
	assign img[40][35] = 1'b0;
	assign img[40][36] = 1'b0;
	assign img[40][37] = 1'b0;
	assign img[40][38] = 1'b0;
	assign img[40][39] = 1'b0;
	assign img[40][40] = 1'b0;
	assign img[40][41] = 1'b0;
	assign img[40][42] = 1'b0;
	assign img[40][43] = 1'b0;
	assign img[40][44] = 1'b0;
	assign img[40][45] = 1'b0;
	assign img[40][46] = 1'b0;
	assign img[40][47] = 1'b0;
	assign img[40][48] = 1'b0;
	assign img[40][49] = 1'b0;
	assign img[40][50] = 1'b0;
	assign img[40][51] = 1'b0;
	assign img[40][52] = 1'b0;
	assign img[40][53] = 1'b0;
	assign img[40][54] = 1'b0;
	assign img[40][55] = 1'b0;
	assign img[40][56] = 1'b0;
	assign img[40][57] = 1'b0;
	assign img[40][58] = 1'b0;
	assign img[40][59] = 1'b0;
	assign img[40][60] = 1'b0;
	assign img[40][61] = 1'b0;
	assign img[40][62] = 1'b0;
	assign img[40][63] = 1'b0;
	assign img[41][0] = 1'b0;
	assign img[41][1] = 1'b0;
	assign img[41][2] = 1'b0;
	assign img[41][3] = 1'b0;
	assign img[41][4] = 1'b0;
	assign img[41][5] = 1'b0;
	assign img[41][6] = 1'b0;
	assign img[41][7] = 1'b0;
	assign img[41][8] = 1'b0;
	assign img[41][9] = 1'b0;
	assign img[41][10] = 1'b0;
	assign img[41][11] = 1'b0;
	assign img[41][12] = 1'b0;
	assign img[41][13] = 1'b0;
	assign img[41][14] = 1'b0;
	assign img[41][15] = 1'b0;
	assign img[41][16] = 1'b0;
	assign img[41][17] = 1'b0;
	assign img[41][18] = 1'b0;
	assign img[41][19] = 1'b0;
	assign img[41][20] = 1'b0;
	assign img[41][21] = 1'b0;
	assign img[41][22] = 1'b0;
	assign img[41][23] = 1'b0;
	assign img[41][24] = 1'b0;
	assign img[41][25] = 1'b0;
	assign img[41][26] = 1'b0;
	assign img[41][27] = 1'b0;
	assign img[41][28] = 1'b0;
	assign img[41][29] = 1'b0;
	assign img[41][30] = 1'b0;
	assign img[41][31] = 1'b0;
	assign img[41][32] = 1'b0;
	assign img[41][33] = 1'b0;
	assign img[41][34] = 1'b0;
	assign img[41][35] = 1'b0;
	assign img[41][36] = 1'b0;
	assign img[41][37] = 1'b0;
	assign img[41][38] = 1'b0;
	assign img[41][39] = 1'b0;
	assign img[41][40] = 1'b0;
	assign img[41][41] = 1'b0;
	assign img[41][42] = 1'b0;
	assign img[41][43] = 1'b0;
	assign img[41][44] = 1'b0;
	assign img[41][45] = 1'b0;
	assign img[41][46] = 1'b0;
	assign img[41][47] = 1'b0;
	assign img[41][48] = 1'b0;
	assign img[41][49] = 1'b0;
	assign img[41][50] = 1'b0;
	assign img[41][51] = 1'b0;
	assign img[41][52] = 1'b0;
	assign img[41][53] = 1'b0;
	assign img[41][54] = 1'b0;
	assign img[41][55] = 1'b0;
	assign img[41][56] = 1'b0;
	assign img[41][57] = 1'b0;
	assign img[41][58] = 1'b0;
	assign img[41][59] = 1'b0;
	assign img[41][60] = 1'b0;
	assign img[41][61] = 1'b1;
	assign img[41][62] = 1'b0;
	assign img[41][63] = 1'b0;
	assign img[42][0] = 1'b0;
	assign img[42][1] = 1'b0;
	assign img[42][2] = 1'b0;
	assign img[42][3] = 1'b0;
	assign img[42][4] = 1'b0;
	assign img[42][5] = 1'b0;
	assign img[42][6] = 1'b0;
	assign img[42][7] = 1'b0;
	assign img[42][8] = 1'b0;
	assign img[42][9] = 1'b0;
	assign img[42][10] = 1'b0;
	assign img[42][11] = 1'b0;
	assign img[42][12] = 1'b0;
	assign img[42][13] = 1'b0;
	assign img[42][14] = 1'b0;
	assign img[42][15] = 1'b0;
	assign img[42][16] = 1'b0;
	assign img[42][17] = 1'b0;
	assign img[42][18] = 1'b0;
	assign img[42][19] = 1'b0;
	assign img[42][20] = 1'b0;
	assign img[42][21] = 1'b0;
	assign img[42][22] = 1'b0;
	assign img[42][23] = 1'b0;
	assign img[42][24] = 1'b0;
	assign img[42][25] = 1'b0;
	assign img[42][26] = 1'b0;
	assign img[42][27] = 1'b0;
	assign img[42][28] = 1'b0;
	assign img[42][29] = 1'b0;
	assign img[42][30] = 1'b0;
	assign img[42][31] = 1'b0;
	assign img[42][32] = 1'b0;
	assign img[42][33] = 1'b0;
	assign img[42][34] = 1'b0;
	assign img[42][35] = 1'b0;
	assign img[42][36] = 1'b0;
	assign img[42][37] = 1'b0;
	assign img[42][38] = 1'b0;
	assign img[42][39] = 1'b0;
	assign img[42][40] = 1'b0;
	assign img[42][41] = 1'b0;
	assign img[42][42] = 1'b0;
	assign img[42][43] = 1'b0;
	assign img[42][44] = 1'b0;
	assign img[42][45] = 1'b0;
	assign img[42][46] = 1'b0;
	assign img[42][47] = 1'b0;
	assign img[42][48] = 1'b0;
	assign img[42][49] = 1'b0;
	assign img[42][50] = 1'b0;
	assign img[42][51] = 1'b0;
	assign img[42][52] = 1'b0;
	assign img[42][53] = 1'b0;
	assign img[42][54] = 1'b0;
	assign img[42][55] = 1'b0;
	assign img[42][56] = 1'b0;
	assign img[42][57] = 1'b0;
	assign img[42][58] = 1'b0;
	assign img[42][59] = 1'b0;
	assign img[42][60] = 1'b0;
	assign img[42][61] = 1'b0;
	assign img[42][62] = 1'b0;
	assign img[42][63] = 1'b0;
	assign img[43][0] = 1'b0;
	assign img[43][1] = 1'b0;
	assign img[43][2] = 1'b0;
	assign img[43][3] = 1'b0;
	assign img[43][4] = 1'b0;
	assign img[43][5] = 1'b0;
	assign img[43][6] = 1'b0;
	assign img[43][7] = 1'b0;
	assign img[43][8] = 1'b0;
	assign img[43][9] = 1'b0;
	assign img[43][10] = 1'b0;
	assign img[43][11] = 1'b0;
	assign img[43][12] = 1'b0;
	assign img[43][13] = 1'b0;
	assign img[43][14] = 1'b0;
	assign img[43][15] = 1'b0;
	assign img[43][16] = 1'b0;
	assign img[43][17] = 1'b0;
	assign img[43][18] = 1'b0;
	assign img[43][19] = 1'b0;
	assign img[43][20] = 1'b0;
	assign img[43][21] = 1'b0;
	assign img[43][22] = 1'b0;
	assign img[43][23] = 1'b0;
	assign img[43][24] = 1'b0;
	assign img[43][25] = 1'b0;
	assign img[43][26] = 1'b0;
	assign img[43][27] = 1'b0;
	assign img[43][28] = 1'b0;
	assign img[43][29] = 1'b0;
	assign img[43][30] = 1'b0;
	assign img[43][31] = 1'b0;
	assign img[43][32] = 1'b0;
	assign img[43][33] = 1'b0;
	assign img[43][34] = 1'b0;
	assign img[43][35] = 1'b0;
	assign img[43][36] = 1'b0;
	assign img[43][37] = 1'b0;
	assign img[43][38] = 1'b0;
	assign img[43][39] = 1'b0;
	assign img[43][40] = 1'b0;
	assign img[43][41] = 1'b0;
	assign img[43][42] = 1'b0;
	assign img[43][43] = 1'b0;
	assign img[43][44] = 1'b0;
	assign img[43][45] = 1'b0;
	assign img[43][46] = 1'b0;
	assign img[43][47] = 1'b0;
	assign img[43][48] = 1'b0;
	assign img[43][49] = 1'b0;
	assign img[43][50] = 1'b0;
	assign img[43][51] = 1'b0;
	assign img[43][52] = 1'b0;
	assign img[43][53] = 1'b0;
	assign img[43][54] = 1'b0;
	assign img[43][55] = 1'b0;
	assign img[43][56] = 1'b0;
	assign img[43][57] = 1'b0;
	assign img[43][58] = 1'b0;
	assign img[43][59] = 1'b0;
	assign img[43][60] = 1'b0;
	assign img[43][61] = 1'b0;
	assign img[43][62] = 1'b0;
	assign img[43][63] = 1'b0;
	assign img[44][0] = 1'b0;
	assign img[44][1] = 1'b0;
	assign img[44][2] = 1'b0;
	assign img[44][3] = 1'b0;
	assign img[44][4] = 1'b1;
	assign img[44][5] = 1'b0;
	assign img[44][6] = 1'b0;
	assign img[44][7] = 1'b0;
	assign img[44][8] = 1'b0;
	assign img[44][9] = 1'b0;
	assign img[44][10] = 1'b0;
	assign img[44][11] = 1'b0;
	assign img[44][12] = 1'b0;
	assign img[44][13] = 1'b0;
	assign img[44][14] = 1'b0;
	assign img[44][15] = 1'b0;
	assign img[44][16] = 1'b0;
	assign img[44][17] = 1'b0;
	assign img[44][18] = 1'b0;
	assign img[44][19] = 1'b1;
	assign img[44][20] = 1'b0;
	assign img[44][21] = 1'b0;
	assign img[44][22] = 1'b0;
	assign img[44][23] = 1'b0;
	assign img[44][24] = 1'b0;
	assign img[44][25] = 1'b0;
	assign img[44][26] = 1'b0;
	assign img[44][27] = 1'b0;
	assign img[44][28] = 1'b0;
	assign img[44][29] = 1'b0;
	assign img[44][30] = 1'b0;
	assign img[44][31] = 1'b0;
	assign img[44][32] = 1'b0;
	assign img[44][33] = 1'b0;
	assign img[44][34] = 1'b0;
	assign img[44][35] = 1'b0;
	assign img[44][36] = 1'b0;
	assign img[44][37] = 1'b0;
	assign img[44][38] = 1'b1;
	assign img[44][39] = 1'b0;
	assign img[44][40] = 1'b0;
	assign img[44][41] = 1'b0;
	assign img[44][42] = 1'b0;
	assign img[44][43] = 1'b0;
	assign img[44][44] = 1'b0;
	assign img[44][45] = 1'b0;
	assign img[44][46] = 1'b0;
	assign img[44][47] = 1'b0;
	assign img[44][48] = 1'b0;
	assign img[44][49] = 1'b0;
	assign img[44][50] = 1'b0;
	assign img[44][51] = 1'b0;
	assign img[44][52] = 1'b0;
	assign img[44][53] = 1'b0;
	assign img[44][54] = 1'b0;
	assign img[44][55] = 1'b0;
	assign img[44][56] = 1'b0;
	assign img[44][57] = 1'b0;
	assign img[44][58] = 1'b0;
	assign img[44][59] = 1'b0;
	assign img[44][60] = 1'b0;
	assign img[44][61] = 1'b0;
	assign img[44][62] = 1'b0;
	assign img[44][63] = 1'b0;
	assign img[45][0] = 1'b0;
	assign img[45][1] = 1'b0;
	assign img[45][2] = 1'b0;
	assign img[45][3] = 1'b0;
	assign img[45][4] = 1'b0;
	assign img[45][5] = 1'b0;
	assign img[45][6] = 1'b0;
	assign img[45][7] = 1'b0;
	assign img[45][8] = 1'b0;
	assign img[45][9] = 1'b0;
	assign img[45][10] = 1'b0;
	assign img[45][11] = 1'b0;
	assign img[45][12] = 1'b0;
	assign img[45][13] = 1'b0;
	assign img[45][14] = 1'b0;
	assign img[45][15] = 1'b0;
	assign img[45][16] = 1'b0;
	assign img[45][17] = 1'b0;
	assign img[45][18] = 1'b0;
	assign img[45][19] = 1'b0;
	assign img[45][20] = 1'b0;
	assign img[45][21] = 1'b0;
	assign img[45][22] = 1'b0;
	assign img[45][23] = 1'b0;
	assign img[45][24] = 1'b0;
	assign img[45][25] = 1'b0;
	assign img[45][26] = 1'b0;
	assign img[45][27] = 1'b0;
	assign img[45][28] = 1'b0;
	assign img[45][29] = 1'b0;
	assign img[45][30] = 1'b0;
	assign img[45][31] = 1'b0;
	assign img[45][32] = 1'b0;
	assign img[45][33] = 1'b0;
	assign img[45][34] = 1'b0;
	assign img[45][35] = 1'b0;
	assign img[45][36] = 1'b0;
	assign img[45][37] = 1'b0;
	assign img[45][38] = 1'b0;
	assign img[45][39] = 1'b0;
	assign img[45][40] = 1'b0;
	assign img[45][41] = 1'b0;
	assign img[45][42] = 1'b0;
	assign img[45][43] = 1'b0;
	assign img[45][44] = 1'b0;
	assign img[45][45] = 1'b0;
	assign img[45][46] = 1'b0;
	assign img[45][47] = 1'b0;
	assign img[45][48] = 1'b0;
	assign img[45][49] = 1'b0;
	assign img[45][50] = 1'b0;
	assign img[45][51] = 1'b0;
	assign img[45][52] = 1'b0;
	assign img[45][53] = 1'b0;
	assign img[45][54] = 1'b0;
	assign img[45][55] = 1'b0;
	assign img[45][56] = 1'b0;
	assign img[45][57] = 1'b0;
	assign img[45][58] = 1'b0;
	assign img[45][59] = 1'b0;
	assign img[45][60] = 1'b0;
	assign img[45][61] = 1'b0;
	assign img[45][62] = 1'b0;
	assign img[45][63] = 1'b0;
	assign img[46][0] = 1'b0;
	assign img[46][1] = 1'b0;
	assign img[46][2] = 1'b0;
	assign img[46][3] = 1'b0;
	assign img[46][4] = 1'b0;
	assign img[46][5] = 1'b0;
	assign img[46][6] = 1'b0;
	assign img[46][7] = 1'b0;
	assign img[46][8] = 1'b0;
	assign img[46][9] = 1'b0;
	assign img[46][10] = 1'b0;
	assign img[46][11] = 1'b0;
	assign img[46][12] = 1'b0;
	assign img[46][13] = 1'b0;
	assign img[46][14] = 1'b0;
	assign img[46][15] = 1'b0;
	assign img[46][16] = 1'b0;
	assign img[46][17] = 1'b0;
	assign img[46][18] = 1'b0;
	assign img[46][19] = 1'b0;
	assign img[46][20] = 1'b0;
	assign img[46][21] = 1'b0;
	assign img[46][22] = 1'b0;
	assign img[46][23] = 1'b0;
	assign img[46][24] = 1'b0;
	assign img[46][25] = 1'b0;
	assign img[46][26] = 1'b0;
	assign img[46][27] = 1'b0;
	assign img[46][28] = 1'b0;
	assign img[46][29] = 1'b0;
	assign img[46][30] = 1'b0;
	assign img[46][31] = 1'b0;
	assign img[46][32] = 1'b0;
	assign img[46][33] = 1'b0;
	assign img[46][34] = 1'b0;
	assign img[46][35] = 1'b0;
	assign img[46][36] = 1'b0;
	assign img[46][37] = 1'b0;
	assign img[46][38] = 1'b0;
	assign img[46][39] = 1'b0;
	assign img[46][40] = 1'b0;
	assign img[46][41] = 1'b0;
	assign img[46][42] = 1'b0;
	assign img[46][43] = 1'b0;
	assign img[46][44] = 1'b0;
	assign img[46][45] = 1'b0;
	assign img[46][46] = 1'b0;
	assign img[46][47] = 1'b0;
	assign img[46][48] = 1'b0;
	assign img[46][49] = 1'b0;
	assign img[46][50] = 1'b0;
	assign img[46][51] = 1'b0;
	assign img[46][52] = 1'b0;
	assign img[46][53] = 1'b0;
	assign img[46][54] = 1'b0;
	assign img[46][55] = 1'b0;
	assign img[46][56] = 1'b0;
	assign img[46][57] = 1'b0;
	assign img[46][58] = 1'b0;
	assign img[46][59] = 1'b0;
	assign img[46][60] = 1'b0;
	assign img[46][61] = 1'b0;
	assign img[46][62] = 1'b0;
	assign img[46][63] = 1'b0;
	assign img[47][0] = 1'b0;
	assign img[47][1] = 1'b0;
	assign img[47][2] = 1'b0;
	assign img[47][3] = 1'b0;
	assign img[47][4] = 1'b0;
	assign img[47][5] = 1'b0;
	assign img[47][6] = 1'b0;
	assign img[47][7] = 1'b0;
	assign img[47][8] = 1'b0;
	assign img[47][9] = 1'b0;
	assign img[47][10] = 1'b0;
	assign img[47][11] = 1'b0;
	assign img[47][12] = 1'b0;
	assign img[47][13] = 1'b0;
	assign img[47][14] = 1'b0;
	assign img[47][15] = 1'b0;
	assign img[47][16] = 1'b0;
	assign img[47][17] = 1'b0;
	assign img[47][18] = 1'b1;
	assign img[47][19] = 1'b0;
	assign img[47][20] = 1'b0;
	assign img[47][21] = 1'b0;
	assign img[47][22] = 1'b0;
	assign img[47][23] = 1'b0;
	assign img[47][24] = 1'b0;
	assign img[47][25] = 1'b0;
	assign img[47][26] = 1'b0;
	assign img[47][27] = 1'b0;
	assign img[47][28] = 1'b0;
	assign img[47][29] = 1'b0;
	assign img[47][30] = 1'b0;
	assign img[47][31] = 1'b0;
	assign img[47][32] = 1'b0;
	assign img[47][33] = 1'b0;
	assign img[47][34] = 1'b0;
	assign img[47][35] = 1'b0;
	assign img[47][36] = 1'b0;
	assign img[47][37] = 1'b0;
	assign img[47][38] = 1'b0;
	assign img[47][39] = 1'b0;
	assign img[47][40] = 1'b0;
	assign img[47][41] = 1'b0;
	assign img[47][42] = 1'b0;
	assign img[47][43] = 1'b0;
	assign img[47][44] = 1'b0;
	assign img[47][45] = 1'b0;
	assign img[47][46] = 1'b0;
	assign img[47][47] = 1'b0;
	assign img[47][48] = 1'b0;
	assign img[47][49] = 1'b0;
	assign img[47][50] = 1'b0;
	assign img[47][51] = 1'b0;
	assign img[47][52] = 1'b0;
	assign img[47][53] = 1'b0;
	assign img[47][54] = 1'b0;
	assign img[47][55] = 1'b0;
	assign img[47][56] = 1'b0;
	assign img[47][57] = 1'b0;
	assign img[47][58] = 1'b0;
	assign img[47][59] = 1'b0;
	assign img[47][60] = 1'b0;
	assign img[47][61] = 1'b0;
	assign img[47][62] = 1'b0;
	assign img[47][63] = 1'b0;
endmodule