module wing(clk, rst, X, Y, mapR, mapG, mapB);

	parameter xbit = 10, ybit = 9;
	input clk, rst;
	input [xbit-1:0] X;
	input [ybit-1:0] Y;
	output [7:0] mapR, mapG, mapB;
	reg [7:0] mapR, mapG, mapB;

	always @(posedge clk, negedge rst) begin
		if(!rst) begin
			mapR <= 8'd255;
			mapG <= 8'd255;
			mapB <= 8'd255;
		end
		else begin
			case(Y)
				`ybit'd0: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd1: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd2: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd3: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd4: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd5: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd6: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd7: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd8: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd9: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd10: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd250, 8'd239, 8'd211};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd246, 8'd234, 8'd196};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd247, 8'd245, 8'd206};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd238, 8'd235, 8'd182};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd11: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd240, 8'd221, 8'd163};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd228, 8'd206, 8'd123};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd188};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd246, 8'd243, 8'd210};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd245, 8'd237, 8'd188};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd232, 8'd207, 8'd123};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd218, 8'd184, 8'd77};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd12: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd234, 8'd201, 8'd122};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd171, 8'd59};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd128};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd248, 8'd230, 8'd168};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd197};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd125};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd233, 8'd174, 8'd48};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd220, 8'd146, 8'd0};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd13: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd239, 8'd188, 8'd97};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd221, 8'd147, 8'd22};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd248, 8'd188, 8'd68};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd114};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd245, 8'd251, 8'd213};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd181};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd128};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd249, 8'd191, 8'd66};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd242, 8'd160, 8'd14};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd243, 8'd144, 8'd0};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd14: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd188, 8'd95};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd241, 8'd142, 8'd15};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd241, 8'd157, 8'd23};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd248, 8'd191, 8'd62};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd125};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd153};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd254, 8'd241, 8'd196};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd248, 8'd245, 8'd202};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd248, 8'd232, 8'd154};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd252, 8'd221, 8'd105};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd249, 8'd197, 8'd59};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd240, 8'd170, 8'd23};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd15};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd253, 8'd157, 8'd21};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd15: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd99};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd21};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd241, 8'd142, 8'd0};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd242, 8'd214, 8'd45};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd244, 8'd222, 8'd87};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd247, 8'd235, 8'd151};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd203};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd250, 8'd227, 8'd160};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd105};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd251, 8'd204, 8'd56};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd242, 8'd180, 8'd17};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd229, 8'd156, 8'd2};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd233, 8'd151, 8'd23};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd247, 8'd163, 8'd51};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd16: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd238, 8'd190, 8'd114};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd244, 8'd159, 8'd42};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd21};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd249, 8'd149, 8'd1};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd238, 8'd190, 8'd28};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd240, 8'd192, 8'd58};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd243, 8'd199, 8'd104};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd250, 8'd215, 8'd149};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd190};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd223};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd221};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd197};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd250, 8'd203, 8'd121};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd245, 8'd207, 8'd84};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd241, 8'd200, 8'd56};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd64};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd247, 8'd165, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd237, 8'd148, 8'd0};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd25};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd242, 8'd163, 8'd42};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd17: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd246, 8'd204, 8'd130};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd240, 8'd163, 8'd45};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd18};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd252, 8'd155, 8'd0};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd239, 8'd172, 8'd32};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd253, 8'd194, 8'd64};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd94};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd243, 8'd213, 8'd103};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd237, 8'd219, 8'd121};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd246, 8'd237, 8'd162};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd207};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd217};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd248, 8'd230, 8'd156};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd239, 8'd216, 8'd110};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd251, 8'd212, 8'd111};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd250, 8'd212, 8'd85};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd247, 8'd199, 8'd63};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd250, 8'd179, 8'd51};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd244, 8'd157, 8'd16};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd243, 8'd155, 8'd0};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd252, 8'd178, 8'd31};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd250, 8'd183, 8'd78};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd18: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd157};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd235, 8'd172, 8'd58};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd248, 8'd164, 8'd16};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd0};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd244, 8'd151, 8'd32};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd56};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd75};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd247, 8'd220, 8'd71};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd231, 8'd217, 8'd68};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd228, 8'd217, 8'd91};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd244, 8'd223, 8'd140};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd179};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd207};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd251, 8'd230, 8'd175};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd244, 8'd215, 8'd137};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd241, 8'd207, 8'd99};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd242, 8'd205, 8'd73};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd100};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd249, 8'd209, 8'd78};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd244, 8'd184, 8'd60};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd241, 8'd155, 8'd36};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd250, 8'd154, 8'd7};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd0};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd246, 8'd185, 8'd43};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd249, 8'd204, 8'd121};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd19: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd187};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd235, 8'd188, 8'd84};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd239, 8'd167, 8'd21};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd2};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd144, 8'd26};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd248, 8'd155, 8'd34};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd252, 8'd187, 8'd57};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd79};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd251, 8'd230, 8'd75};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd229, 8'd211, 8'd65};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd234, 8'd205, 8'd85};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd254, 8'd216, 8'd119};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd245, 8'd224, 8'd167};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd254, 8'd235, 8'd192};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd224};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd253, 8'd247, 8'd169};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd245, 8'd230, 8'd111};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd236, 8'd209, 8'd80};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd235, 8'd201, 8'd78};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd245, 8'd208, 8'd94};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd109};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd84};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd239, 8'd193, 8'd56};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd235, 8'd162, 8'd47};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd240, 8'd140, 8'd26};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd8};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd5};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd231, 8'd187, 8'd56};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd241, 8'd219, 8'd162};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd20: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd238, 8'd206, 8'd119};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd233, 8'd174, 8'd38};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd6};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd18};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd246, 8'd146, 8'd22};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd239, 8'd161, 8'd52};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd92};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd102};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd86};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd244, 8'd210, 8'd77};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd251, 8'd212, 8'd85};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd228, 8'd210, 8'd84};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd238, 8'd220, 8'd112};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd252, 8'd234, 8'd158};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd203};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd249, 8'd229, 8'd170};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd237, 8'd215, 8'd104};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd233, 8'd208, 8'd63};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd237, 8'd209, 8'd63};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd246, 8'd216, 8'd86};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd251, 8'd223, 8'd113};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd252, 8'd227, 8'd126};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd246, 8'd204, 8'd58};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd229, 8'd173, 8'd34};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd238, 8'd158, 8'd37};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd252, 8'd149, 8'd31};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd16};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd250, 8'd179, 8'd11};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd219, 8'd187, 8'd74};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd245, 8'd236, 8'd203};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd21: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd246, 8'd228, 8'd162};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd62};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd248, 8'd171, 8'd13};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd9};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd24};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd237, 8'd151, 8'd48};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd234, 8'd165, 8'd74};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd251, 8'd197, 8'd101};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd112};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd107};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd94};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd247, 8'd228, 8'd74};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd236, 8'd217, 8'd76};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd232, 8'd211, 8'd94};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd241, 8'd219, 8'd133};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd186};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd234};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd122};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd245, 8'd211, 8'd104};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd240, 8'd207, 8'd92};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd242, 8'd210, 8'd97};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd249, 8'd218, 8'd112};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd253, 8'd224, 8'd120};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd250, 8'd224, 8'd111};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd244, 8'd223, 8'd98};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd231, 8'd171, 8'd38};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd233, 8'd166, 8'd25};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd252, 8'd170, 8'd34};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd40};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd23};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd232, 8'd167, 8'd23};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd225, 8'd200, 8'd110};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd22: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd253, 8'd247, 8'd199};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd235, 8'd192, 8'd88};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd241, 8'd167, 8'd20};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd6};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd23};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd245, 8'd159, 8'd38};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd48};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd240, 8'd175, 8'd71};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd107};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd130};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd135};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd110};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd251, 8'd223, 8'd97};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd238, 8'd210, 8'd84};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd234, 8'd208, 8'd89};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd241, 8'd217, 8'd117};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd249, 8'd231, 8'd157};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd253, 8'd240, 8'd195};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd253, 8'd244, 8'd215};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd197, 8'd210, 8'd216};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd139, 8'd156, 8'd163};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd139, 8'd158, 8'd165};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd152, 8'd181, 8'd185};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd196, 8'd224, 8'd227};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd206, 8'd224, 8'd224};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd196, 8'd221, 8'd218};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd196, 8'd221, 8'd218};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd205, 8'd223, 8'd223};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd253, 8'd245, 8'd209};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd250, 8'd235, 8'd176};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd248, 8'd225, 8'd147};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd128};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd85};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd89};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd248, 8'd221, 8'd106};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd253, 8'd229, 8'd131};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd148};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd135};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd246, 8'd205, 8'd99};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd236, 8'd192, 8'd67};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd239, 8'd155, 8'd43};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd28};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd26};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd36};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd244, 8'd161, 8'd33};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd232, 8'd175, 8'd59};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd250, 8'd227, 8'd160};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd23: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd236, 8'd197, 8'd102};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd236, 8'd163, 8'd25};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd251, 8'd176, 8'd5};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd253, 8'd175, 8'd17};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd254, 8'd169, 8'd27};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd248, 8'd165, 8'd35};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd241, 8'd173, 8'd50};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd239, 8'd192, 8'd86};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd242, 8'd215, 8'd134};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd245, 8'd230, 8'd171};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd248, 8'd213, 8'd131};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd125};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd110};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd92};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd243, 8'd217, 8'd81};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd232, 8'd213, 8'd93};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd233, 8'd221, 8'd123};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd239, 8'd231, 8'd148};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd169, 8'd188, 8'd194};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd143, 8'd166, 8'd172};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd166, 8'd193, 8'd200};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd139, 8'd179, 8'd181};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd123, 8'd158, 8'd160};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd149, 8'd179, 8'd181};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd217, 8'd237, 8'd238};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd219, 8'd230, 8'd232};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd139, 8'd161, 8'd159};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd138, 8'd167, 8'd163};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd137, 8'd166, 8'd162};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd138, 8'd160, 8'd158};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd217, 8'd228, 8'd230};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd251, 8'd248, 8'd213};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd247, 8'd238, 8'd179};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd241, 8'd223, 8'd137};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd237, 8'd209, 8'd99};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd234, 8'd200, 8'd76};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd118};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd104};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd238, 8'd222, 8'd101};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd249, 8'd237, 8'd125};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd150};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd141};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd245, 8'd189, 8'd94};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd222, 8'd153, 8'd50};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd60};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd33};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd253, 8'd174, 8'd9};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd251, 8'd171, 8'd24};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd239, 8'd163, 8'd43};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd248, 8'd194, 8'd96};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd199};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd24: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd253, 8'd230, 8'd189};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd221, 8'd190, 8'd136};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd36};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd249, 8'd177, 8'd13};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd242, 8'd177, 8'd23};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd250, 8'd168, 8'd56};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd52};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd250, 8'd161, 8'd31};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd242, 8'd183, 8'd67};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd239, 8'd205, 8'd133};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd174};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd247, 8'd225, 8'd152};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd242, 8'd215, 8'd136};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd131};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd121};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd252, 8'd222, 8'd98};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd236, 8'd213, 8'd73};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd228, 8'd208, 8'd59};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd239, 8'd217, 8'd131};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd247, 8'd227, 8'd154};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd186};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd193, 8'd221, 8'd222};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd150, 8'd173, 8'd187};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd171, 8'd206};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd119, 8'd105, 8'd154};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd145, 8'd159, 8'd206};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd136, 8'd162, 8'd195};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd108, 8'd146, 8'd157};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd147, 8'd181, 8'd180};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd189, 8'd199, 8'd209};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd127, 8'd134, 8'd153};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd148, 8'd159, 8'd189};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd160, 8'd184, 8'd218};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd150, 8'd187, 8'd213};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd148, 8'd186, 8'd199};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd148, 8'd172, 8'd174};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd211};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd188};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd248, 8'd232, 8'd144};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd232, 8'd209, 8'd95};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd231, 8'd201, 8'd77};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd243, 8'd213, 8'd93};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd253, 8'd222, 8'd114};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd252, 8'd224, 8'd125};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd157};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd244, 8'd227, 8'd149};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd245, 8'd229, 8'd154};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd160};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd136};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd240, 8'd185, 8'd85};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd241, 8'd163, 8'd52};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd44};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd235, 8'd181, 8'd21};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd247, 8'd165, 8'd37};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd40};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd22};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd225, 8'd181, 8'd58};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd244, 8'd224, 8'd173};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd25: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd253, 8'd237, 8'd203};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd228, 8'd205, 8'd161};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd246, 8'd170, 8'd50};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd252, 8'd182, 8'd26};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd21};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd254, 8'd170, 8'd38};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd159, 8'd41};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd251, 8'd166, 8'd37};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd245, 8'd178, 8'd61};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd240, 8'd185, 8'd102};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd246, 8'd230, 8'd152};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd161};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd161};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd251, 8'd226, 8'd146};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd247, 8'd220, 8'd129};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd223, 8'd117};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd102};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd251, 8'd218, 8'd85};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd245, 8'd212, 8'd83};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd244, 8'd215, 8'd97};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd246, 8'd222, 8'd126};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd254, 8'd236, 8'd170};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd159, 8'd183, 8'd187};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd154, 8'd172, 8'd192};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd158, 8'd157, 8'd197};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd134, 8'd115, 8'd170};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd154, 8'd119, 8'd187};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd136, 8'd124, 8'd174};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd152, 8'd164, 8'd190};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd143, 8'd163, 8'd170};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd208, 8'd219, 8'd215};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd138, 8'd155, 8'd163};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd160, 8'd164, 8'd189};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd141, 8'd133, 8'd180};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd121, 8'd118, 8'd173};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd89, 8'd101, 8'd149};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd171, 8'd195, 8'd223};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd125, 8'd148, 8'd154};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd246, 8'd229, 8'd160};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd239, 8'd218, 8'd137};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd236, 8'd211, 8'd108};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd246, 8'd216, 8'd96};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd101};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd112};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd253, 8'd224, 8'd122};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd245, 8'd219, 8'd126};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd243, 8'd225, 8'd149};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd168};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd167};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd248, 8'd212, 8'd136};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd231, 8'd184, 8'd96};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd236, 8'd171, 8'd67};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd250, 8'd171, 8'd50};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd39};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd250, 8'd180, 8'd33};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd28};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd251, 8'd166, 8'd15};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd237, 8'd170, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd239, 8'd203, 8'd115};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd253, 8'd239, 8'd212};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd26: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd239, 8'd228, 8'd198};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd235, 8'd181, 8'd91};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd245, 8'd182, 8'd43};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd9};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd16};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd33};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd246, 8'd167, 8'd36};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd246, 8'd167, 8'd48};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd250, 8'd167, 8'd65};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd228, 8'd201, 8'd110};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd248, 8'd226, 8'd143};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd171};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd173};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd246, 8'd225, 8'd158};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd249, 8'd222, 8'd141};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd128};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd117};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd85};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd82};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd242, 8'd210, 8'd89};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd239, 8'd216, 8'd112};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd242, 8'd229, 8'd150};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd250, 8'd242, 8'd193};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd163, 8'd177, 8'd186};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd179, 8'd189, 8'd216};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd104, 8'd94, 8'd144};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd156, 8'd130, 8'd193};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd181, 8'd98, 8'd186};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd114, 8'd63, 8'd132};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd165, 8'd153, 8'd193};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd140, 8'd152, 8'd166};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd179, 8'd190, 8'd186};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd145, 8'd173, 8'd177};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd138, 8'd137, 8'd169};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd106, 8'd75, 8'd143};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd182, 8'd139, 8'd228};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd147, 8'd123, 8'd201};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd165, 8'd167, 8'd216};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd170, 8'd194, 8'd206};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd153, 8'd186, 8'd175};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd206};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd231, 8'd162};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd133};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd247, 8'd209, 8'd112};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd236, 8'd199, 8'd93};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd237, 8'd202, 8'd84};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd99};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd118};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd127};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd250, 8'd226, 8'd136};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd247, 8'd224, 8'd146};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd245, 8'd227, 8'd155};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd168};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd153};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd241, 8'd182, 8'd102};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd227, 8'd157, 8'd62};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd242, 8'd162, 8'd49};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd42};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd31};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd38};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd15};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd240, 8'd172, 8'd1};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd228, 8'd183, 8'd68};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd252, 8'd231, 8'd186};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd27: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd243, 8'd214, 8'd158};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd236, 8'd184, 8'd72};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd247, 8'd168, 8'd3};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd4};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd240, 8'd166, 8'd35};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd245, 8'd155, 8'd33};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd37};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd227, 8'd167, 8'd69};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd234, 8'd184, 8'd99};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd247, 8'd212, 8'd144};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd183};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd188};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd246, 8'd228, 8'd164};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd245, 8'd222, 8'd142};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd254, 8'd227, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd134};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd124};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd251, 8'd219, 8'd106};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd240, 8'd215, 8'd89};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd233, 8'd212, 8'd87};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd237, 8'd217, 8'd104};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd248, 8'd230, 8'd132};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd153};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd169, 8'd177, 8'd190};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd173, 8'd178, 8'd208};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd118, 8'd105, 8'd158};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd144, 8'd115, 8'd181};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd164, 8'd84, 8'd173};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd47, 8'd117};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd159, 8'd154, 8'd194};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd130, 8'd149, 8'd166};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd181, 8'd192, 8'd188};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd143, 8'd181, 8'd182};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd117, 8'd115, 8'd152};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd94, 8'd47, 8'd127};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd195, 8'd128, 8'd234};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd148, 8'd96, 8'd196};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd118, 8'd104, 8'd165};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd182, 8'd205, 8'd221};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd138, 8'd180, 8'd166};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd187};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd251, 8'd224, 8'd143};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd243, 8'd213, 8'd103};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd238, 8'd204, 8'd78};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd95};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd252, 8'd211, 8'd93};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd250, 8'd218, 8'd99};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd254, 8'd229, 8'd113};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd252, 8'd233, 8'd128};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd247, 8'd232, 8'd141};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd248, 8'd234, 8'd159};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd176};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd164};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd248, 8'd210, 8'd139};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd243, 8'd181, 8'd106};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd245, 8'd163, 8'd77};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd252, 8'd160, 8'd57};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd40};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd254, 8'd172, 8'd28};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd251, 8'd177, 8'd20};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd21};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd9};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd239, 8'd189, 8'd40};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd237, 8'd210, 8'd139};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd28: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd252, 8'd242, 8'd215};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd239, 8'd201, 8'd126};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd240, 8'd172, 8'd35};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd252, 8'd176, 8'd5};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd25};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd246, 8'd172, 8'd41};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd252, 8'd158, 8'd32};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd16};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd249, 8'd153, 8'd50};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd239, 8'd156, 8'd64};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd104};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd252, 8'd212, 8'd153};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd182};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd252, 8'd240, 8'd180};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd236, 8'd162};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd238, 8'd233, 8'd151};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd239, 8'd219, 8'd156};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd147};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd127};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd254, 8'd229, 8'd102};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd79};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd247, 8'd210, 8'd69};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd249, 8'd205, 8'd70};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd253, 8'd205, 8'd77};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd231, 8'd220, 8'd141};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd243, 8'd232, 8'd168};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd206};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd170, 8'd177, 8'd187};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd141, 8'd147, 8'd173};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd181, 8'd172, 8'd217};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd128, 8'd104, 8'd164};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd103, 8'd68, 8'd134};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd98, 8'd90, 8'd141};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd159, 8'd184, 8'd214};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd111, 8'd149, 8'd160};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd214};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd110, 8'd154, 8'd153};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd153, 8'd158, 8'd190};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd101, 8'd59, 8'd133};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd124, 8'd59, 8'd159};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd128, 8'd77, 8'd170};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd162, 8'd147, 8'd204};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd131, 8'd150, 8'd165};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd160, 8'd201, 8'd187};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd205};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd248, 8'd233, 8'd166};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd243, 8'd223, 8'd128};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd241, 8'd216, 8'd100};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd244, 8'd213, 8'd86};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd213, 8'd83};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd253, 8'd214, 8'd85};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd105};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd116};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd125};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd246, 8'd232, 8'd135};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd242, 8'd235, 8'd147};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd249, 8'd241, 8'd168};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd254, 8'd243, 8'd179};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd183};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd141};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd233, 8'd180, 8'd100};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd229, 8'd153, 8'd67};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd252, 8'd158, 8'd58};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd55};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd38};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd253, 8'd171, 8'd23};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd248, 8'd175, 8'd18};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd253, 8'd163, 8'd7};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd242, 8'd176, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd119};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd253, 8'd241, 8'd215};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd29: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd251, 8'd231, 8'd196};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd245, 8'd200, 8'd107};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd235, 8'd177, 8'd31};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd243, 8'd174, 8'd21};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd50};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd43};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd6};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd46};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd55};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd244, 8'd161, 8'd69};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd236, 8'd173, 8'd94};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd247, 8'd205, 8'd133};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd167};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd174};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd241, 8'd239, 8'd164};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd238, 8'd234, 8'd147};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd236, 8'd230, 8'd136};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd241, 8'd227, 8'd120};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd249, 8'd227, 8'd108};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd103};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd98};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd89};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd82};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd231, 8'd207, 8'd101};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd233, 8'd209, 8'd113};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd238, 8'd217, 8'd138};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd251, 8'd232, 8'd176};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd213};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd224, 8'd234, 8'd236};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd160, 8'd172, 8'd186};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd137, 8'd140, 8'd171};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd156, 8'd147, 8'd190};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd90, 8'd104, 8'd141};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd90, 8'd121, 8'd149};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd138, 8'd186, 8'd200};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd108, 8'd153, 8'd159};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd224, 8'd235, 8'd231};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd110, 8'd156, 8'd154};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd166, 8'd182, 8'd205};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd87, 8'd70, 8'd122};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd112, 8'd81, 8'd149};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd180, 8'd158, 8'd220};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd168, 8'd168, 8'd206};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd139, 8'd156, 8'd166};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd198, 8'd221, 8'd213};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd191, 8'd191, 8'd191};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd244, 8'd223, 8'd170};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd242, 8'd220, 8'd145};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd240, 8'd216, 8'd108};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd240, 8'd214, 8'd77};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd244, 8'd214, 8'd66};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd250, 8'd217, 8'd76};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd96};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd111};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd254, 8'd223, 8'd117};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd253, 8'd229, 8'd129};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd247, 8'd232, 8'd141};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd241, 8'd235, 8'd151};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd252, 8'd244, 8'd169};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd179};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd166};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd243, 8'd210, 8'd143};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd241, 8'd179, 8'd94};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd238, 8'd167, 8'd75};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd245, 8'd159, 8'd56};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd44};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd39};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd35};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd254, 8'd176, 8'd28};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd245, 8'd174, 8'd24};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd243, 8'd172, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd237, 8'd189, 8'd89};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd196};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd30: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd252, 8'd234, 8'd188};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd235, 8'd196, 8'd79};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd239, 8'd172, 8'd31};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd48};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd47};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd244, 8'd174, 8'd14};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd43};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd45};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd250, 8'd161, 8'd43};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd236, 8'd153, 8'd49};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd238, 8'd167, 8'd75};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd252, 8'd199, 8'd119};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd155};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd168};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd254, 8'd241, 8'd149};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd248, 8'd233, 8'd142};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd245, 8'd224, 8'd133};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd247, 8'd221, 8'd128};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd126};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd124};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd116};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd110};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd100};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd93};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd237, 8'd204, 8'd89};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd236, 8'd209, 8'd102};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd243, 8'd222, 8'd131};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd253, 8'd236, 8'd167};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd198};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd214};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd210, 8'd231, 8'd232};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd115, 8'd133, 8'd147};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd152, 8'd160, 8'd183};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd121, 8'd157, 8'd173};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd82, 8'd126, 8'd137};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd126, 8'd173, 8'd179};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd113, 8'd148, 8'd154};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd217, 8'd228, 8'd224};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd112, 8'd158, 8'd156};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd146, 8'd176, 8'd186};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd74, 8'd89, 8'd110};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd132, 8'd144, 8'd170};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd149, 8'd167, 8'd189};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd107, 8'd126, 8'd140};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd207, 8'd218, 8'd222};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd195, 8'd201, 8'd199};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd131, 8'd131, 8'd131};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd187};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd252, 8'd227, 8'd160};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd248, 8'd223, 8'd143};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd237, 8'd208, 8'd106};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd242, 8'd210, 8'd99};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd248, 8'd212, 8'd90};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd253, 8'd216, 8'd84};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd88};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd101};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd254, 8'd223, 8'd115};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd253, 8'd224, 8'd124};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd128};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd250, 8'd226, 8'd136};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd245, 8'd230, 8'd147};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd249, 8'd235, 8'd160};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd162};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd146};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd250, 8'd196, 8'd110};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd236, 8'd171, 8'd81};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd244, 8'd157, 8'd60};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd252, 8'd165, 8'd59};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd49};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd33};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd254, 8'd169, 8'd26};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd251, 8'd176, 8'd35};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd244, 8'd171, 8'd33};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd239, 8'd190, 8'd85};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd251, 8'd222, 8'd166};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd31: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd247, 8'd218, 8'd124};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd245, 8'd177, 8'd42};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd38};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd254, 8'd176, 8'd42};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd244, 8'd191, 8'd27};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd243, 8'd186, 8'd37};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd245, 8'd174, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd246, 8'd163, 8'd25};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd247, 8'd153, 8'd31};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd239, 8'd146, 8'd42};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd234, 8'd156, 8'd71};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd250, 8'd190, 8'd120};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd164};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd159};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd164};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd169};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd161};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd145};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd245, 8'd219, 8'd126};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd244, 8'd220, 8'd112};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd246, 8'd223, 8'd107};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd101};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd93};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd79};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd240, 8'd212, 8'd69};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd230, 8'd208, 8'd73};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd229, 8'd212, 8'd98};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd237, 8'd221, 8'd133};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd245, 8'd231, 8'd158};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd88, 8'd108, 8'd119};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd133, 8'd168, 8'd174};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd95, 8'd134, 8'd139};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd156, 8'd191, 8'd195};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd115, 8'd135, 8'd142};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd197, 8'd201, 8'd210};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd201, 8'd212, 8'd208};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd101, 8'd145, 8'd144};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd146, 8'd184, 8'd185};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd77, 8'd115, 8'd116};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd126, 8'd168, 8'd166};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd85, 8'd130, 8'd125};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd170, 8'd205, 8'd199};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd197, 8'd203, 8'd201};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd130, 8'd136, 8'd134};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd89};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd212};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd177};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd246, 8'd220, 8'd135};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd238, 8'd208, 8'd94};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd232, 8'd202, 8'd70};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd82};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd86};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd94};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd102};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd113};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd122};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd248, 8'd222, 8'd127};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd246, 8'd226, 8'd131};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd138};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd254, 8'd228, 8'd143};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd252, 8'd233, 8'd154};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd161};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd140};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd239, 8'd185, 8'd95};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd235, 8'd157, 8'd57};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd239, 8'd147, 8'd38};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd55};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd47};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd35};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd253, 8'd171, 8'd25};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd249, 8'd174, 8'd23};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd248, 8'd173, 8'd28};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd244, 8'd170, 8'd35};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd243, 8'd168, 8'd40};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd241, 8'd207, 8'd135};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd219};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd32: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd232, 8'd211, 8'd156};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd229, 8'd180, 8'd85};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd248, 8'd170, 8'd34};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd13};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd223, 8'd186, 8'd0};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd232, 8'd173, 8'd17};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd252, 8'd163, 8'd43};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd53};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd40};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd249, 8'd156, 8'd35};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd61};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd237, 8'd174, 8'd94};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd127};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd134};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd246, 8'd224, 8'd141};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd239, 8'd227, 8'd145};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd239, 8'd224, 8'd139};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd248, 8'd219, 8'd127};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd117};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd110};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd94};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd92};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd251, 8'd211, 8'd89};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd245, 8'd209, 8'd86};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd244, 8'd209, 8'd83};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd246, 8'd208, 8'd83};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd248, 8'd209, 8'd82};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd252, 8'd208, 8'd83};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd243, 8'd217, 8'd133};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd251, 8'd227, 8'd157};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd194};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd169, 8'd173, 8'd184};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd167, 8'd173, 8'd189};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd221, 8'd227, 8'd249};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd162, 8'd164, 8'd163};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd97, 8'd136, 8'd135};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd147, 8'd181, 8'd182};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd134, 8'd158, 8'd162};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd95, 8'd108, 8'd116};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd120, 8'd127, 8'd133};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd133, 8'd143, 8'd144};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd123, 8'd148, 8'd153};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd155, 8'd188, 8'd193};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd132, 8'd169, 8'd175};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd121, 8'd150, 8'd158};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd154, 8'd166, 8'd178};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd190, 8'd200, 8'd201};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd146, 8'd157, 8'd159};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd127, 8'd141, 8'd144};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd107, 8'd126, 8'd107};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd210};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd187};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd225, 8'd149};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd240, 8'd210, 8'd112};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd237, 8'd204, 8'd88};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd242, 8'd207, 8'd81};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd249, 8'd214, 8'd84};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd254, 8'd221, 8'd88};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd96};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd213, 8'd96};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd246, 8'd215, 8'd99};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd247, 8'd221, 8'd110};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd251, 8'd226, 8'd123};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd130};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd135};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd133};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd245, 8'd222, 8'd155};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd165};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd161};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd124};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd251, 8'd179, 8'd71};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd240, 8'd160, 8'd37};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd249, 8'd161, 8'd38};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd55};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd247, 8'd161, 8'd26};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd250, 8'd162, 8'd38};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd251, 8'd168, 8'd38};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd248, 8'd174, 8'd13};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd241, 8'd181, 8'd0};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd239, 8'd183, 8'd10};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd240, 8'd184, 8'd75};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd245, 8'd183, 8'd134};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd33: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd199};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd254, 8'd215, 8'd140};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd247, 8'd183, 8'd73};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd242, 8'd161, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd247, 8'd183, 8'd0};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd253, 8'd181, 8'd17};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd38};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd249, 8'd163, 8'd44};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd252, 8'd163, 8'd47};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd50};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd49};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd239, 8'd154, 8'd45};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd239, 8'd168, 8'd76};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd248, 8'd187, 8'd98};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd125};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd143};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd143};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd249, 8'd225, 8'd129};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd248, 8'd219, 8'd117};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd109};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd103};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd100};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd251, 8'd216, 8'd96};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd93};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd247, 8'd216, 8'd91};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd251, 8'd216, 8'd90};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd89};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd90};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd243, 8'd216, 8'd99};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd236, 8'd212, 8'd106};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd231, 8'd209, 8'd123};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd236, 8'd218, 8'd154};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd248, 8'd237, 8'd191};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd172, 8'd180, 8'd182};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd115, 8'd124, 8'd129};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd170, 8'd183, 8'd191};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd212, 8'd225, 8'd234};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd182, 8'd184, 8'd183};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd84, 8'd113, 8'd108};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd100, 8'd122, 8'd120};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd91, 8'd105, 8'd106};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd71, 8'd74, 8'd79};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd80, 8'd79, 8'd84};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd213, 8'd217, 8'd218};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd83};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd88, 8'd102, 8'd105};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd107, 8'd131, 8'd133};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd119, 8'd150, 8'd152};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd93, 8'd118, 8'd123};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd188, 8'd197, 8'd206};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd185, 8'd195, 8'd197};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd158, 8'd169, 8'd173};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd157, 8'd172, 8'd179};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd107, 8'd122, 8'd129};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd126, 8'd132, 8'd146};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd237, 8'd217, 8'd131};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd238, 8'd215, 8'd122};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd241, 8'd210, 8'd104};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd243, 8'd206, 8'd91};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd246, 8'd204, 8'd83};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd251, 8'd207, 8'd84};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd253, 8'd211, 8'd91};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd96};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd200, 8'd85};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd96};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd108};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd254, 8'd227, 8'd114};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd247, 8'd225, 8'd116};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd246, 8'd223, 8'd121};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd251, 8'd227, 8'd129};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd137};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd138};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd251, 8'd206, 8'd125};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd236, 8'd179, 8'd98};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd230, 8'd161, 8'd66};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd235, 8'd157, 8'd46};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd247, 8'd161, 8'd40};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd51};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd62};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd242, 8'd170, 8'd36};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd245, 8'd164, 8'd29};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd21};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd9};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd251, 8'd177, 8'd4};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd235, 8'd179, 8'd40};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd239, 8'd202, 8'd124};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd204};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd34: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd198};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd249, 8'd206, 8'd137};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd232, 8'd176, 8'd91};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd250, 8'd164, 8'd3};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd17};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd32};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd247, 8'd178, 8'd39};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd244, 8'd168, 8'd48};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd251, 8'd164, 8'd48};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd31};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd14};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd245, 8'd153, 8'd44};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd245, 8'd158, 8'd53};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd250, 8'd171, 8'd76};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd104};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd125};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd131};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd243, 8'd226, 8'd120};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd227, 8'd219, 8'd108};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd248, 8'd211, 8'd104};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd105};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd220, 8'd107};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd108};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd104};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd97};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd254, 8'd216, 8'd89};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd253, 8'd212, 8'd86};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd76};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd243, 8'd214, 8'd74};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd236, 8'd207, 8'd77};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd229, 8'd202, 8'd89};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd230, 8'd205, 8'd112};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd239, 8'd215, 8'd145};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd178};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd199};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd201};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd84, 8'd99, 8'd94};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd139, 8'd158, 8'd152};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd164, 8'd185, 8'd178};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd220, 8'd224, 8'd227};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd213, 8'd215, 8'd214};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd87, 8'd99, 8'd89};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd46, 8'd51, 8'd44};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd47, 8'd42, 8'd38};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd42, 8'd30, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd27, 8'd13, 8'd13};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd185, 8'd175, 8'd176};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd179, 8'd175, 8'd174};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd25, 8'd19, 8'd19};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd77, 8'd73, 8'd72};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd76, 8'd85, 8'd82};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd90, 8'd109, 8'd107};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd103, 8'd119, 8'd119};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd205, 8'd214, 8'd219};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd136, 8'd149, 8'd157};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd145, 8'd159, 8'd170};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd153, 8'd169, 8'd182};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd77, 8'd95, 8'd107};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd167, 8'd166, 8'd180};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd252, 8'd249, 8'd198};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd240, 8'd230, 8'd158};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd228, 8'd211, 8'd123};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd222, 8'd199, 8'd105};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd232, 8'd197, 8'd69};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd239, 8'd202, 8'd70};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd248, 8'd208, 8'd74};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd79};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd87};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd94};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd101};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd107};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd97};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd96};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd251, 8'd214, 8'd99};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd104};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd249, 8'd221, 8'd111};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd250, 8'd223, 8'd116};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd223, 8'd118};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd250, 8'd223, 8'd120};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd254, 8'd196, 8'd88};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd238, 8'd173, 8'd73};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd224, 8'd150, 8'd53};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd228, 8'd145, 8'd39};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd247, 8'd158, 8'd38};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd43};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd49};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd253, 8'd158, 8'd52};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd230, 8'd167, 8'd26};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd253, 8'd178, 8'd27};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd15};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd254, 8'd164, 8'd6};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd250, 8'd173, 8'd43};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd125};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd209};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd35: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd203};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd250, 8'd221, 8'd181};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd240, 8'd167, 8'd54};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd241, 8'd170, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd12};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd20};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd35};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd162, 8'd37};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd25};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd17};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd41};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd251, 8'd159, 8'd36};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd241, 8'd146, 8'd36};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd240, 8'd152, 8'd52};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd248, 8'd174, 8'd79};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd254, 8'd200, 8'd102};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd114};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd243, 8'd225, 8'd117};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd251, 8'd214, 8'd110};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd250, 8'd216, 8'd109};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd250, 8'd218, 8'd107};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd250, 8'd221, 8'd104};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd100};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd94};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd251, 8'd213, 8'd88};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd84};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd84};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd79};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd252, 8'd214, 8'd71};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd241, 8'd202, 8'd63};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd230, 8'd189, 8'd63};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd227, 8'd183, 8'd76};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd233, 8'd185, 8'd100};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd240, 8'd190, 8'd117};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd245, 8'd219, 8'd168};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd202};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd86, 8'd105, 8'd103};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd133, 8'd154, 8'd147};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd140, 8'd163, 8'd153};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd171, 8'd180, 8'd189};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd224, 8'd231, 8'd239};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd142, 8'd138, 8'd126};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd53, 8'd40, 8'd31};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd62, 8'd37, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd59, 8'd28, 8'd25};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd26, 8'd0, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd121, 8'd101, 8'd100};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd126, 8'd110, 8'd110};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd17, 8'd0, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd29, 8'd4, 8'd0};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd29, 8'd18, 8'd12};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd12, 8'd17, 8'd10};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd140, 8'd146, 8'd142};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd214, 8'd219, 8'd223};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd147, 8'd157, 8'd166};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd143, 8'd159, 8'd172};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd161, 8'd179, 8'd193};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd125, 8'd143, 8'd157};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd65, 8'd83, 8'd97};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd198, 8'd205, 8'd189};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd250, 8'd236, 8'd201};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd239, 8'd220, 8'd152};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd226, 8'd202, 8'd106};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd222, 8'd189, 8'd76};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd227, 8'd187, 8'd66};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd234, 8'd188, 8'd66};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd241, 8'd198, 8'd60};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd247, 8'd204, 8'd65};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd74};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd82};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd91};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd97};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd252, 8'd212, 8'd98};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd247, 8'd206, 8'd98};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd102};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd253, 8'd221, 8'd100};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd251, 8'd216, 8'd98};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd253, 8'd216, 8'd101};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd103};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd100};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd247, 8'd196, 8'd91};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd238, 8'd185, 8'd81};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd238, 8'd156, 8'd48};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd241, 8'd154, 8'd51};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd248, 8'd155, 8'd52};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd47};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd37};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd28};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd248, 8'd159, 8'd31};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd238, 8'd165, 8'd10};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd249, 8'd177, 8'd17};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd248, 8'd177, 8'd25};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd241, 8'd176, 8'd56};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd251, 8'd201, 8'd130};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd216};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd36: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd249, 8'd212, 8'd159};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd232, 8'd187, 8'd86};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd227, 8'd166, 8'd15};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd247, 8'd165, 8'd0};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd14};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd33};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd33};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd246, 8'd171, 8'd26};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd252, 8'd180, 8'd33};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd35};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd253, 8'd161, 8'd36};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd243, 8'd145, 8'd34};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd235, 8'd139, 8'd37};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd237, 8'd155, 8'd56};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd185, 8'd85};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd109};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd115};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd111};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd213, 8'd105};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd247, 8'd211, 8'd97};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd93};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd249, 8'd213, 8'd91};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd254, 8'd216, 8'd93};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd93};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd109};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd92};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd246, 8'd196, 8'd71};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd244, 8'd191, 8'd59};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd244, 8'd190, 8'd56};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd242, 8'd182, 8'd58};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd235, 8'd172, 8'd59};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd227, 8'd162, 8'd58};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd208, 8'd170, 8'd59};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd223, 8'd192, 8'd99};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd240, 8'd221, 8'd152};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd248, 8'd239, 8'd196};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd90, 8'd107, 8'd114};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd115, 8'd136, 8'd139};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd137, 8'd162, 8'd159};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd149, 8'd161, 8'd173};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd176, 8'd189, 8'd198};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd198, 8'd184, 8'd173};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd83, 8'd56, 8'd47};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd90, 8'd49, 8'd43};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd89, 8'd40, 8'd35};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd51, 8'd6, 8'd3};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd47, 8'd17, 8'd15};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd239, 8'd229, 8'd227};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd239, 8'd221, 8'd219};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd69, 8'd43, 8'd42};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd42, 8'd8, 8'd7};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd94, 8'd47, 8'd39};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd97, 8'd69, 8'd58};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd45, 8'd38, 8'd28};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd172, 8'd181, 8'd188};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd131, 8'd148, 8'd158};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd172, 8'd191, 8'd205};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd162, 8'd181, 8'd195};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd100, 8'd116, 8'd129};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd86, 8'd100, 8'd111};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd215, 8'd226, 8'd212};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd187};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd248, 8'd209, 8'd152};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd225, 8'd182, 8'd103};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd213, 8'd166, 8'd62};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd218, 8'd164, 8'd42};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd232, 8'd171, 8'd44};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd244, 8'd179, 8'd53};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd251, 8'd183, 8'd60};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd242, 8'd192, 8'd77};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd244, 8'd197, 8'd79};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd205, 8'd84};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd212, 8'd87};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd248, 8'd214, 8'd88};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd243, 8'd214, 8'd88};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd239, 8'd209, 8'd85};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd235, 8'd207, 8'd84};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd238, 8'd220, 8'd92};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd249, 8'd225, 8'd99};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd106};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd102};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd86};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd248, 8'd174, 8'd67};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd241, 8'd158, 8'd54};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd240, 8'd151, 8'd49};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd245, 8'd147, 8'd46};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd252, 8'd152, 8'd54};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd59};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd46};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd23};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd11};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd11};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd250, 8'd173, 8'd19};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd13};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd233, 8'd165, 8'd20};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd229, 8'd183, 8'd71};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd248, 8'd225, 8'd158};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd231};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd37: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd248, 8'd231, 8'd177};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd241, 8'd194, 8'd90};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd23};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd248, 8'd159, 8'd7};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd24};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd252, 8'd176, 8'd38};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd235, 8'd171, 8'd37};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd240, 8'd174, 8'd26};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd250, 8'd175, 8'd32};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd38};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd39};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd250, 8'd148, 8'd37};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd247, 8'd146, 8'd42};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd154, 8'd52};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd65};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd84};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd90};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd98};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd103};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd103};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd100};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd93};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd251, 8'd209, 8'd89};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd116};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd105};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd247, 8'd193, 8'd87};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd241, 8'd184, 8'd69};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd238, 8'd178, 8'd58};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd236, 8'd172, 8'd49};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd233, 8'd167, 8'd45};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd233, 8'd164, 8'd43};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd225, 8'd173, 8'd35};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd209, 8'd159, 8'd34};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd200, 8'd153, 8'd49};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd211, 8'd170, 8'd88};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd238, 8'd203, 8'd137};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd174};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd183};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd179};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd133};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd91, 8'd110, 8'd117};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd153, 8'd174, 8'd179};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd155, 8'd174, 8'd181};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd139, 8'd156, 8'd163};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd183, 8'd196, 8'd202};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd227, 8'd209, 8'd205};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd107, 8'd76, 8'd73};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd98, 8'd47, 8'd44};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd108, 8'd44, 8'd42};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd77, 8'd18, 8'd14};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd28, 8'd0, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd184, 8'd169, 8'd164};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd183, 8'd159, 8'd155};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd41, 8'd3, 8'd0};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd66, 8'd20, 8'd20};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd96, 8'd33, 8'd26};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd102, 8'd59, 8'd50};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd85, 8'd68, 8'd58};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd185, 8'd193, 8'd195};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd153, 8'd168, 8'd175};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd163, 8'd183, 8'd194};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd178, 8'd200, 8'd211};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd132, 8'd151, 8'd158};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd92, 8'd106, 8'd109};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd129, 8'd137, 8'd139};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd251, 8'd243, 8'd196};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd245, 8'd229, 8'd167};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd232, 8'd209, 8'd133};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd234, 8'd206, 8'd123};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd219, 8'd160, 8'd66};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd220, 8'd158, 8'd59};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd223, 8'd157, 8'd47};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd229, 8'd158, 8'd40};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd237, 8'd163, 8'd42};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd48};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd246, 8'd170, 8'd58};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd248, 8'd171, 8'd63};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd240, 8'd186, 8'd88};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd241, 8'd192, 8'd90};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd243, 8'd201, 8'd93};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd245, 8'd209, 8'd95};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd246, 8'd216, 8'd94};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd247, 8'd218, 8'd92};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd247, 8'd218, 8'd90};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd246, 8'd217, 8'd87};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd222, 8'd97};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd92};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd252, 8'd200, 8'd82};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd252, 8'd182, 8'd68};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd56};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd249, 8'd152, 8'd45};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd251, 8'd146, 8'd41};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd251, 8'd144, 8'd38};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd252, 8'd157, 8'd49};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd253, 8'd156, 8'd51};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd254, 8'd158, 8'd48};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd36};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd20};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd252, 8'd175, 8'd9};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd244, 8'd175, 8'd10};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd239, 8'd173, 8'd16};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd248, 8'd174, 8'd43};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd241, 8'd188, 8'd84};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd242, 8'd222, 8'd161};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd248, 8'd255, 8'd233};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd38: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd252, 8'd246, 8'd214};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd235, 8'd226, 8'd183};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd244, 8'd232, 8'd180};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd197};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd196};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd249, 8'd204, 8'd121};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd239, 8'd179, 8'd55};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd243, 8'd172, 8'd28};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd248, 8'd173, 8'd28};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd249, 8'd172, 8'd34};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd32};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd248, 8'd164, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd251, 8'd162, 8'd32};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd38};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd45};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd44};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd253, 8'd147, 8'd37};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd243, 8'd136, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd237, 8'd149, 8'd39};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd245, 8'd163, 8'd53};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd71};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd89};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd98};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd99};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd94};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd248, 8'd203, 8'd88};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd252, 8'd204, 8'd94};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd254, 8'd203, 8'd96};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd251, 8'd198, 8'd96};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd241, 8'd183, 8'd83};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd229, 8'd167, 8'd66};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd223, 8'd159, 8'd53};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd226, 8'd160, 8'd48};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd232, 8'd165, 8'd50};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd229, 8'd160, 8'd41};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd228, 8'd155, 8'd40};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd223, 8'd145, 8'd36};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd215, 8'd136, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd211, 8'd137, 8'd38};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd219, 8'd159, 8'd61};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd238, 8'd192, 8'd96};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd254, 8'd218, 8'd122};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd183};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd250, 8'd244, 8'd186};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd160, 8'd171, 8'd173};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd78, 8'd93, 8'd96};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd146, 8'd166, 8'd165};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd160, 8'd184, 8'd188};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd142, 8'd163, 8'd166};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd155, 8'd173, 8'd175};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd204, 8'd218, 8'd219};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd146, 8'd114, 8'd117};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd104, 8'd48, 8'd49};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd133, 8'd61, 8'd62};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd102, 8'd34, 8'd31};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd42, 8'd0, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd126, 8'd107, 8'd101};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd99, 8'd72, 8'd65};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd49, 8'd4, 8'd1};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd83, 8'd27, 8'd26};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd124, 8'd49, 8'd43};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd101, 8'd51, 8'd42};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd150, 8'd130, 8'd119};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd203};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd157, 8'd173, 8'd173};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd156, 8'd177, 8'd182};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd174, 8'd201, 8'd210};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd165, 8'd190, 8'd197};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd106, 8'd124, 8'd126};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd93, 8'd99, 8'd95};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd166, 8'd168, 8'd157};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd249, 8'd233, 8'd197};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd175};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd239, 8'd212, 8'd123};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd238, 8'd198, 8'd87};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd217, 8'd166, 8'd38};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd209, 8'd150, 8'd14};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd206, 8'd133, 8'd18};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd215, 8'd139, 8'd27};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd225, 8'd144, 8'd36};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd227, 8'd146, 8'd39};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd226, 8'd147, 8'd44};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd228, 8'd155, 8'd53};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd237, 8'd169, 8'd70};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd245, 8'd181, 8'd83};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd241, 8'd178, 8'd73};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd244, 8'd186, 8'd79};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd249, 8'd198, 8'd89};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd253, 8'd210, 8'd97};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd100};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd98};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd93};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd89};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd85};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd253, 8'd180, 8'd69};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd241, 8'd156, 8'd47};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd239, 8'd144, 8'd36};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd245, 8'd145, 8'd34};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd253, 8'd151, 8'd40};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd42};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd42};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd29};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd249, 8'd164, 8'd35};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd38};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd251, 8'd169, 8'd33};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd251, 8'd175, 8'd27};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd248, 8'd179, 8'd26};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd241, 8'd179, 8'd34};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd236, 8'd176, 8'd43};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd239, 8'd201, 8'd120};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd183};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd247, 8'd230, 8'd176};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd243, 8'd221, 8'd163};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd176};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd39: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd241, 8'd232, 8'd173};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd210, 8'd199, 8'd119};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd216, 8'd204, 8'd106};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd245, 8'd233, 8'd125};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd210};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd128};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd245, 8'd189, 8'd50};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd248, 8'd168, 8'd17};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd17};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd36};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd35};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd253, 8'd159, 8'd33};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd251, 8'd162, 8'd34};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd254, 8'd162, 8'd35};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd36};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd36};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd35};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd234, 8'd133, 8'd19};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd234, 8'd140, 8'd26};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd236, 8'd152, 8'd38};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd239, 8'd170, 8'd53};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd245, 8'd186, 8'd70};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd251, 8'd200, 8'd85};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd97};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd102};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd243, 8'd201, 8'd63};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd239, 8'd194, 8'd67};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd235, 8'd185, 8'd74};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd233, 8'd179, 8'd83};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd234, 8'd175, 8'd85};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd233, 8'd170, 8'd77};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd227, 8'd163, 8'd63};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd221, 8'd158, 8'd52};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd221, 8'd141, 8'd52};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd232, 8'd143, 8'd49};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd239, 8'd140, 8'd38};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd236, 8'd130, 8'd20};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd226, 8'd127, 8'd10};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd220, 8'd140, 8'd17};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd227, 8'd169, 8'd43};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd234, 8'd194, 8'd63};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd243, 8'd235, 8'd136};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd231, 8'd225, 8'd139};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd242, 8'd238, 8'd175};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd246, 8'd244, 8'd206};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd205};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd71, 8'd86, 8'd79};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd118, 8'd137, 8'd131};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd153, 8'd179, 8'd178};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd163, 8'd187, 8'd187};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd156, 8'd176, 8'd177};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd169, 8'd183, 8'd184};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd216, 8'd226, 8'd228};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd166, 8'd133, 8'd142};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd96, 8'd37, 8'd43};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd137, 8'd63, 8'd64};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd101, 8'd30, 8'd28};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd70, 8'd19, 8'd15};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd70, 8'd50, 8'd43};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd216, 8'd216, 8'd208};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd231, 8'd221, 8'd212};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd34, 8'd3, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd70, 8'd21, 8'd17};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd92, 8'd31, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd158, 8'd77, 8'd73};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd102, 8'd47, 8'd40};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd195, 8'd171, 8'd161};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd164, 8'd179, 8'd176};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd163, 8'd183, 8'd182};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd163, 8'd188, 8'd193};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd159, 8'd188, 8'd194};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd154, 8'd179, 8'd183};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd102, 8'd118, 8'd115};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd90, 8'd93, 8'd82};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd182, 8'd179, 8'd162};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd239, 8'd216, 8'd162};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd234, 8'd210, 8'd148};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd236, 8'd210, 8'd133};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd249, 8'd214, 8'd120};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd238, 8'd190, 8'd79};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd246, 8'd182, 8'd58};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd228, 8'd147, 8'd12};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd215, 8'd125, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd219, 8'd142, 8'd26};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd218, 8'd137, 8'd29};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd218, 8'd134, 8'd36};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd222, 8'd138, 8'd48};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd225, 8'd149, 8'd63};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd225, 8'd159, 8'd72};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd220, 8'd165, 8'd74};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd215, 8'd166, 8'd71};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd237, 8'd167, 8'd46};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd242, 8'd176, 8'd56};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd249, 8'd190, 8'd72};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd254, 8'd201, 8'd85};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd90};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd254, 8'd201, 8'd87};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd251, 8'd194, 8'd81};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd248, 8'd186, 8'd75};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd247, 8'd140, 8'd42};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd251, 8'd143, 8'd44};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd144, 8'd44};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd40};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd252, 8'd146, 8'd36};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd248, 8'd151, 8'd36};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd249, 8'd161, 8'd38};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd250, 8'd168, 8'd43};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd249, 8'd180, 8'd14};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd253, 8'd180, 8'd25};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd253, 8'd178, 8'd35};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd248, 8'd173, 8'd32};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd242, 8'd171, 8'd27};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd240, 8'd177, 8'd38};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd247, 8'd187, 8'd65};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd254, 8'd196, 8'd89};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd253, 8'd248, 8'd208};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd253, 8'd240, 8'd188};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd164};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd237, 8'd206, 8'd126};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd230, 8'd194, 8'd108};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd253, 8'd213, 8'd125};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd40: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd190};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd217, 8'd169, 8'd45};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd241, 8'd178, 8'd15};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd252, 8'd197, 8'd34};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd251, 8'd199, 8'd77};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd127};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd193};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd176};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd244, 8'd201, 8'd86};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd235, 8'd189, 8'd18};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd242, 8'd168, 8'd7};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd244, 8'd176, 8'd17};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd245, 8'd180, 8'd26};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd241, 8'd176, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd238, 8'd167, 8'd27};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd243, 8'd161, 8'd26};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd34};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd41};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd45};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd39};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd146, 8'd28};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd238, 8'd138, 8'd18};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd230, 8'd137, 8'd18};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd234, 8'd153, 8'd38};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd252, 8'd180, 8'd72};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd97};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd251, 8'd200, 8'd73};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd238, 8'd178, 8'd58};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd242, 8'd176, 8'd63};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd235, 8'd175, 8'd61};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd232, 8'd183, 8'd65};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd212, 8'd166, 8'd46};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd219, 8'd160, 8'd40};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd220, 8'd148, 8'd28};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd219, 8'd144, 8'd43};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd218, 8'd140, 8'd42};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd219, 8'd135, 8'd39};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd218, 8'd129, 8'd35};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd212, 8'd122, 8'd25};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd213, 8'd126, 8'd21};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd235, 8'd151, 8'd37};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd59};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd252, 8'd196, 8'd75};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd102};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd122};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd238, 8'd200, 8'd125};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd173};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd241, 8'd220, 8'd177};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd99, 8'd101, 8'd80};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd95, 8'd115, 8'd113};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd146, 8'd172, 8'd171};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd160, 8'd186, 8'd187};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd166, 8'd189, 8'd195};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd149, 8'd169, 8'd178};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd160, 8'd174, 8'd183};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd211, 8'd192, 8'd188};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd69, 8'd30, 8'd25};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd122, 8'd69, 8'd63};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd94, 8'd37, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd73, 8'd26, 8'd20};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd36, 8'd5, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd165, 8'd144, 8'd139};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd157, 8'd138, 8'd131};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd41, 8'd7, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd74, 8'd27, 8'd19};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd88, 8'd33, 8'd26};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd125, 8'd73, 8'd62};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd85, 8'd51, 8'd41};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd217, 8'd227, 8'd228};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd158, 8'd170, 8'd168};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd167, 8'd182, 8'd177};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd157, 8'd178, 8'd171};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd164, 8'd190, 8'd187};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd167, 8'd192, 8'd199};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd130, 8'd146, 8'd161};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd96, 8'd95, 8'd100};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd129, 8'd113, 8'd90};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd193, 8'd169, 8'd123};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd227, 8'd189, 8'd127};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd220, 8'd179, 8'd99};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd240, 8'd196, 8'd87};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd75};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd243, 8'd177, 8'd39};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd244, 8'd164, 8'd39};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd218, 8'd125, 8'd22};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd225, 8'd124, 8'd36};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd219, 8'd131, 8'd41};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd220, 8'd132, 8'd42};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd219, 8'd134, 8'd41};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd218, 8'd138, 8'd43};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd216, 8'd142, 8'd45};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd217, 8'd149, 8'd48};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd219, 8'd157, 8'd54};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd220, 8'd163, 8'd58};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd223, 8'd179, 8'd48};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd217, 8'd169, 8'd41};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd225, 8'd171, 8'd47};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd249, 8'd187, 8'd68};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd80};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd69};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd241, 8'd145, 8'd43};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd227, 8'd125, 8'd27};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd127, 8'd34};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd247, 8'd136, 8'd29};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd244, 8'd150, 8'd24};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd244, 8'd168, 8'd23};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd250, 8'd178, 8'd32};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd254, 8'd176, 8'd40};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd251, 8'd165, 8'd44};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd250, 8'd155, 8'd47};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd245, 8'd167, 8'd31};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd27};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd243, 8'd171, 8'd25};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd228, 8'd170, 8'd45};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd225, 8'd188, 8'd99};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd240, 8'd225, 8'd170};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd223};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd216};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd159};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd245, 8'd217, 8'd92};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd244, 8'd195, 8'd56};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd48};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd254, 8'd187, 8'd21};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd229, 8'd174, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd112};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd41: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd189};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd219, 8'd168, 8'd43};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd242, 8'd173, 8'd10};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd253, 8'd190, 8'd27};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd238, 8'd195, 8'd56};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd241, 8'd200, 8'd84};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd246, 8'd209, 8'd120};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd250, 8'd221, 8'd153};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd254, 8'd235, 8'd177};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd204};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd222};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd254, 8'd229, 8'd173};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd242, 8'd214, 8'd130};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd236, 8'd173, 8'd57};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd242, 8'd174, 8'd49};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd250, 8'd172, 8'd36};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd27};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd24};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd254, 8'd163, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd247, 8'd161, 8'd38};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd244, 8'd160, 8'd46};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd60};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd53};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd250, 8'd149, 8'd43};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd244, 8'd142, 8'd32};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd240, 8'd138, 8'd28};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd238, 8'd140, 8'd29};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd238, 8'd143, 8'd33};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd237, 8'd147, 8'd37};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd248, 8'd179, 8'd60};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd250, 8'd174, 8'd62};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd66};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd229, 8'd157, 8'd49};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd223, 8'd163, 8'd51};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd216, 8'd159, 8'd44};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd229, 8'd159, 8'd45};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd224, 8'd143, 8'd28};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd211, 8'd131, 8'd32};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd212, 8'd129, 8'd33};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd215, 8'd128, 8'd33};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd214, 8'd123, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd205, 8'd115, 8'd18};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd206, 8'd119, 8'd14};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd226, 8'd144, 8'd32};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd251, 8'd172, 8'd54};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd237, 8'd175, 8'd42};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd248, 8'd193, 8'd74};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd253, 8'd209, 8'd104};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd234, 8'd193, 8'd103};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd235, 8'd197, 8'd122};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd220, 8'd198, 8'd141};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd115, 8'd114, 8'd83};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd83, 8'd101, 8'd87};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd117, 8'd141, 8'd145};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd166, 8'd189, 8'd195};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd184, 8'd207, 8'd215};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd158, 8'd178, 8'd187};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd156, 8'd170, 8'd179};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd196, 8'd203, 8'd209};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd107, 8'd70, 8'd62};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd129, 8'd76, 8'd68};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd114, 8'd57, 8'd48};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd97, 8'd47, 8'd38};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd43, 8'd6, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd88, 8'd59, 8'd55};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd104, 8'd79, 8'd74};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd45, 8'd6, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd75, 8'd22, 8'd16};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd101, 8'd40, 8'd35};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd118, 8'd68, 8'd61};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd119, 8'd86, 8'd79};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd188, 8'd198, 8'd200};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd167, 8'd181, 8'd184};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd172, 8'd188, 8'd185};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd176, 8'd199, 8'd193};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd175, 8'd204, 8'd200};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd153, 8'd180, 8'd187};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd112, 8'd128, 8'd141};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd94, 8'd92, 8'd93};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd129, 8'd109, 8'd84};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd178, 8'd148, 8'd98};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd205, 8'd158, 8'd88};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd220, 8'd173, 8'd85};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd232, 8'd180, 8'd68};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd230, 8'd172, 8'd39};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd242, 8'd174, 8'd39};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd231, 8'd151, 8'd28};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd207, 8'd115, 8'd14};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd205, 8'd107, 8'd20};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd209, 8'd117, 8'd16};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd212, 8'd123, 8'd23};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd219, 8'd131, 8'd31};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd224, 8'd138, 8'd37};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd222, 8'd143, 8'd40};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd220, 8'd146, 8'd41};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd219, 8'd148, 8'd42};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd217, 8'd150, 8'd43};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd244, 8'd173, 8'd57};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd243, 8'd170, 8'd55};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd169, 8'd58};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd248, 8'd163, 8'd54};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd239, 8'd146, 8'd40};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd230, 8'd129, 8'd25};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd236, 8'd128, 8'd29};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd249, 8'd137, 8'd39};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd45};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd49};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd49};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd253, 8'd163, 8'd41};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd245, 8'd160, 8'd31};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd243, 8'd160, 8'd22};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd247, 8'd164, 8'd22};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd27};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd22};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd246, 8'd169, 8'd15};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd230, 8'd161, 8'd21};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd232, 8'd177, 8'd58};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd247, 8'd210, 8'd122};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd191};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd249, 8'd242, 8'd198};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd240, 8'd228, 8'd178};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd246, 8'd226, 8'd153};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd230, 8'd211, 8'd93};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd240, 8'd210, 8'd62};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd54};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd32};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd238, 8'd166, 8'd4};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd225, 8'd169, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd252, 8'd210, 8'd112};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd42: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd187};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd225, 8'd167, 8'd44};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd244, 8'd164, 8'd5};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd252, 8'd178, 8'd17};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd247, 8'd206, 8'd52};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd249, 8'd201, 8'd55};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd253, 8'd197, 8'd60};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd67};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd86};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd126};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd252, 8'd231, 8'd174};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd250, 8'd239, 8'd211};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd150};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd252, 8'd201, 8'd109};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd246, 8'd171, 8'd52};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd251, 8'd160, 8'd17};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd10};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd22};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd253, 8'd178, 8'd35};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd238, 8'd174, 8'd40};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd247, 8'd167, 8'd54};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd243, 8'd158, 8'd49};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd243, 8'd147, 8'd44};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd247, 8'd144, 8'd43};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd143, 8'd41};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd254, 8'd139, 8'd32};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd244, 8'd130, 8'd16};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd235, 8'd122, 8'd4};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd212, 8'd119, 8'd13};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd230, 8'd131, 8'd29};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd251, 8'd149, 8'd51};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd239, 8'd147, 8'd48};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd238, 8'd161, 8'd57};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd228, 8'd154, 8'd47};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd229, 8'd147, 8'd39};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd222, 8'd127, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd209, 8'd122, 8'd25};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd210, 8'd122, 8'd25};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd213, 8'd120, 8'd27};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd209, 8'd116, 8'd23};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd200, 8'd107, 8'd12};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd199, 8'd112, 8'd9};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd221, 8'd139, 8'd29};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd247, 8'd170, 8'd54};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd243, 8'd170, 8'd29};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd236, 8'd171, 8'd41};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd236, 8'd183, 8'd67};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd230, 8'd181, 8'd78};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd208, 8'd164, 8'd75};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd202, 8'd173, 8'd103};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd136, 8'd129, 8'd85};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd81, 8'd93, 8'd69};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd91, 8'd111, 8'd120};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd162, 8'd182, 8'd191};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd189, 8'd211, 8'd222};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd170, 8'd190, 8'd199};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd158, 8'd175, 8'd182};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd166, 8'd177, 8'd179};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd200, 8'd204, 8'd203};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd140, 8'd108, 8'd97};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd107, 8'd58, 8'd44};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd112, 8'd54, 8'd42};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd97, 8'd40, 8'd29};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd52, 8'd5, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd38, 8'd0, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd214, 8'd205, 8'd198};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd214, 8'd196, 8'd192};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd67, 8'd36, 8'd31};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd80, 8'd32, 8'd28};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd100, 8'd41, 8'd37};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd134, 8'd66, 8'd63};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd106, 8'd58, 8'd58};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd166, 8'd137, 8'd133};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd202, 8'd200, 8'd201};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd171, 8'd182, 8'd188};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd175, 8'd193, 8'd203};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd174, 8'd194, 8'd192};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd188, 8'd215, 8'd208};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd178, 8'd209, 8'd204};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd132, 8'd161, 8'd165};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd95, 8'd109, 8'd118};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd102, 8'd94, 8'd91};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd138, 8'd109, 8'd79};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd166, 8'd125, 8'd71};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd195, 8'd137, 8'd55};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd225, 8'd165, 8'd69};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd227, 8'd166, 8'd51};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd223, 8'd156, 8'd26};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd253, 8'd180, 8'd51};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd216, 8'd135, 8'd18};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd198, 8'd108, 8'd11};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd202, 8'd107, 8'd23};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd224, 8'd127, 8'd20};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd215, 8'd118, 8'd13};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd205, 8'd110, 8'd4};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd205, 8'd114, 8'd9};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd216, 8'd128, 8'd22};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd228, 8'd143, 8'd37};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd236, 8'd151, 8'd45};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd236, 8'd153, 8'd49};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd254, 8'd150, 8'd55};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd243, 8'd136, 8'd40};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd233, 8'd125, 8'd27};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd234, 8'd122, 8'd24};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd236, 8'd122, 8'd23};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd242, 8'd124, 8'd24};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd253, 8'd136, 8'd33};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd148, 8'd44};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd50};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd48};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd45};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd43};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd36};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd27};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd18};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd249, 8'd178, 8'd12};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd241, 8'd168, 8'd4};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd239, 8'd174, 8'd32};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd241, 8'd193, 8'd85};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd153};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd218};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd204};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd246, 8'd228, 8'd156};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd239, 8'd216, 8'd110};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd234, 8'd209, 8'd82};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd238, 8'd215, 8'd83};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd222, 8'd198, 8'd38};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd248, 8'd209, 8'd43};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd49};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd247, 8'd167, 8'd16};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd234, 8'd160, 8'd0};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd231, 8'd175, 8'd40};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd244, 8'd203, 8'd111};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd43: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd188};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd231, 8'd171, 8'd51};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd246, 8'd159, 8'd2};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd251, 8'd168, 8'd10};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd41};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd47};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd50};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd45};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd247, 8'd201, 8'd46};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd240, 8'd202, 8'd65};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd238, 8'd207, 8'd99};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd237, 8'd211, 8'd127};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd157};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd182};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd218};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd172};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd243, 8'd207, 8'd113};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd237, 8'd181, 8'd60};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd239, 8'd171, 8'd24};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd245, 8'd173, 8'd9};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd180, 8'd7};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd253, 8'd183, 8'd7};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd249, 8'd172, 8'd32};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd246, 8'd162, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd247, 8'd153, 8'd31};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd253, 8'd149, 8'd36};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd41};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd35};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd254, 8'd139, 8'd22};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd246, 8'd131, 8'd12};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd227, 8'd113, 8'd16};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd222, 8'd103, 8'd9};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd225, 8'd106, 8'd16};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd222, 8'd114, 8'd23};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd232, 8'd142, 8'd45};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd134, 8'd32};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd220, 8'd128, 8'd25};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd229, 8'd127, 8'd26};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd219, 8'd129, 8'd32};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd219, 8'd126, 8'd31};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd218, 8'd123, 8'd31};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd212, 8'd114, 8'd25};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd196, 8'd101, 8'd9};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd189, 8'd99, 8'd2};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd204, 8'd121, 8'd15};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd225, 8'd147, 8'd36};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd47};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd238, 8'd160, 8'd34};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd213, 8'd146, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd222, 8'd160, 8'd57};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd206, 8'd149, 8'd59};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd195, 8'd152, 8'd83};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd149, 8'd130, 8'd88};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd102, 8'd101, 8'd80};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd86, 8'd102, 8'd115};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd136, 8'd154, 8'd166};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd173, 8'd193, 8'd204};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd180, 8'd200, 8'd209};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd173, 8'd192, 8'd198};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd164, 8'd180, 8'd180};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd176, 8'd187, 8'd181};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd206, 8'd213, 8'd205};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd180, 8'd152, 8'd140};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd91, 8'd45, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd111, 8'd55, 8'd40};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd87, 8'd29, 8'd17};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd68, 8'd15, 8'd7};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd52, 8'd3, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd146, 8'd135, 8'd129};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd136, 8'd112, 8'd108};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd33, 8'd0, 8'd0};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd79, 8'd28, 8'd24};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd95, 8'd32, 8'd27};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd124, 8'd55, 8'd50};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd92, 8'd50, 8'd52};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd205, 8'd181, 8'd179};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd194, 8'd179, 8'd172};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd174, 8'd170, 8'd171};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd179, 8'd192, 8'd200};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd176, 8'd198, 8'd212};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd178, 8'd198, 8'd197};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd183, 8'd210, 8'd205};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd158, 8'd190, 8'd185};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd111, 8'd139, 8'd142};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd90, 8'd101, 8'd105};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd115, 8'd98, 8'd90};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd150, 8'd107, 8'd72};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd164, 8'd108, 8'd49};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd198, 8'd123, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd219, 8'd146, 8'd44};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd222, 8'd147, 8'd32};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd238, 8'd163, 8'd38};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd46};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd197, 8'd111, 8'd2};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd192, 8'd101, 8'd8};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd210, 8'd115, 8'd33};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd221, 8'd114, 8'd16};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd218, 8'd116, 8'd16};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd215, 8'd117, 8'd16};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd215, 8'd121, 8'd21};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd218, 8'd126, 8'd25};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd224, 8'd132, 8'd33};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd229, 8'd135, 8'd37};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd232, 8'd138, 8'd40};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd245, 8'd123, 8'd38};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd223, 8'd101, 8'd15};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd213, 8'd89, 8'd0};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd226, 8'd103, 8'd9};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd250, 8'd128, 8'd29};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd39};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd40};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd39};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd45};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd33};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd23};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd20};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd27};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd33};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd247, 8'd178, 8'd38};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd236, 8'd177, 8'd37};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd246, 8'd194, 8'd84};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd253, 8'd213, 8'd125};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd185};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd215};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd210};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd192};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd247, 8'd230, 8'd161};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd238, 8'd215, 8'd122};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd236, 8'd205, 8'd88};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd244, 8'd205, 8'd65};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd252, 8'd209, 8'd53};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd245, 8'd212, 8'd59};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd248, 8'd211, 8'd45};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd51};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd254, 8'd177, 8'd39};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd247, 8'd158, 8'd14};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd250, 8'd174, 8'd13};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd241, 8'd187, 8'd52};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd242, 8'd205, 8'd116};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd44: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd195};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd238, 8'd178, 8'd64};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd247, 8'd159, 8'd7};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd249, 8'd164, 8'd9};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd244, 8'd163, 8'd9};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd251, 8'd180, 8'd38};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd253, 8'd200, 8'd68};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd247, 8'd213, 8'd77};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd238, 8'd214, 8'd66};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd235, 8'd210, 8'd55};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd243, 8'd209, 8'd58};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd252, 8'd209, 8'd68};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd81};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd242, 8'd209, 8'd102};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd241, 8'd213, 8'd139};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd243, 8'd225, 8'd179};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd241, 8'd234, 8'd179};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd227, 8'd201, 8'd114};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd223, 8'd174, 8'd53};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd237, 8'd166, 8'd14};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd254, 8'd167, 8'd0};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd12};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd15};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd18};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd28};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd253, 8'd151, 8'd27};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd244, 8'd145, 8'd25};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd237, 8'd141, 8'd21};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd249, 8'd125, 8'd29};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd237, 8'd108, 8'd16};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd228, 8'd100, 8'd11};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd224, 8'd111, 8'd19};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd244, 8'd152, 8'd53};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd221, 8'd140, 8'd35};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd204, 8'd117, 8'd11};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd201, 8'd104, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd213, 8'd124, 8'd24};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd215, 8'd120, 8'd26};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd218, 8'd120, 8'd29};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd216, 8'd116, 8'd28};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd202, 8'd104, 8'd15};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd186, 8'd91, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd184, 8'd96, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd193, 8'd108, 8'd2};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd50};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd249, 8'd158, 8'd51};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd205, 8'd126, 8'd25};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd205, 8'd129, 8'd35};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd197, 8'd125, 8'd41};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd183, 8'd123, 8'd61};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd152, 8'd114, 8'd78};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd127, 8'd108, 8'd94};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd89, 8'd102, 8'd111};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd105, 8'd122, 8'd132};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd153, 8'd171, 8'd183};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd188, 8'd208, 8'd217};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd183, 8'd204, 8'd209};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd171, 8'd191, 8'd190};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd169, 8'd186, 8'd180};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd165, 8'd178, 8'd169};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd217, 8'd217, 8'd191};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd232, 8'd210, 8'd199};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd105, 8'd66, 8'd51};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd128, 8'd76, 8'd62};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd103, 8'd47, 8'd34};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd83, 8'd29, 8'd19};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd64, 8'd14, 8'd7};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd85, 8'd74, 8'd68};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd245, 8'd231, 8'd228};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd51, 8'd26, 8'd22};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd30, 8'd0, 8'd0};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd80, 8'd30, 8'd23};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd107, 8'd48, 8'd40};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd130, 8'd67, 8'd58};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd96, 8'd60, 8'd60};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd231};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd245, 8'd234, 8'd214};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd240, 8'd225, 8'd206};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd217, 8'd201, 8'd188};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd159};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd171, 8'd172, 8'd174};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd184, 8'd198, 8'd207};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd176, 8'd198, 8'd211};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd190, 8'd209, 8'd213};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd169, 8'd195, 8'd194};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd132, 8'd163, 8'd158};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd98, 8'd124, 8'd123};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd94, 8'd98, 8'd99};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd120, 8'd92, 8'd80};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd149, 8'd91, 8'd51};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd166, 8'd88, 8'd24};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd190, 8'd103, 8'd6};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd212, 8'd125, 8'd22};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd220, 8'd134, 8'd23};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd246, 8'd159, 8'd44};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd216, 8'd126, 8'd16};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd183, 8'd91, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd190, 8'd95, 8'd5};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd203, 8'd106, 8'd25};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd216, 8'd106, 8'd21};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd218, 8'd112, 8'd26};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd215, 8'd117, 8'd28};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd204, 8'd113, 8'd20};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd197, 8'd110, 8'd15};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd204, 8'd117, 8'd20};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd227, 8'd137, 8'd41};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd248, 8'd155, 8'd60};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd236, 8'd118, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd227, 8'd108, 8'd18};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd226, 8'd105, 8'd12};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd237, 8'd118, 8'd18};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd246, 8'd131, 8'd24};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd246, 8'd141, 8'd24};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd247, 8'd151, 8'd28};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd252, 8'd163, 8'd35};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd252, 8'd175, 8'd33};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd24};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd10};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd3};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd248, 8'd169, 8'd14};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd242, 8'd175, 8'd45};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd241, 8'd187, 8'd89};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd245, 8'd198, 8'd120};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd198};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd222};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd212};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd192};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd252, 8'd233, 8'd157};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd239, 8'd222, 8'd130};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd228, 8'd211, 8'd95};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd226, 8'd207, 8'd68};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd236, 8'd211, 8'd59};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd253, 8'd216, 8'd66};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd77};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd84};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd80};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd73};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd59};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd240, 8'd151, 8'd33};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd21};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd19};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd235, 8'd187, 8'd53};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd248, 8'd220, 8'd137};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd45: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd253, 8'd248, 8'd208};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd243, 8'd191, 8'd82};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd246, 8'd164, 8'd16};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd246, 8'd167, 8'd14};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd242, 8'd148, 8'd0};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd246, 8'd165, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd247, 8'd191, 8'd78};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd244, 8'd212, 8'd103};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd240, 8'd220, 8'd95};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd242, 8'd220, 8'd74};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd250, 8'd216, 8'd56};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd50};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd250, 8'd203, 8'd73};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd248, 8'd204, 8'd81};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd245, 8'd206, 8'd87};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd92};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd241, 8'd220, 8'd105};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd246, 8'd230, 8'd135};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd181};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd215};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd249, 8'd243, 8'd227};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd169};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd189, 8'd109};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd72};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd241, 8'd165, 8'd19};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd246, 8'd166, 8'd17};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd169, 8'd15};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd16};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd20};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd26};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd240, 8'd152, 8'd28};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd232, 8'd145, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd237, 8'd115, 8'd14};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd244, 8'd117, 8'd20};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd239, 8'd116, 8'd22};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd232, 8'd128, 8'd31};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd80};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd252, 8'd185, 8'd72};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd219, 8'd148, 8'd32};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd192, 8'd112, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd189, 8'd103, 8'd2};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd189, 8'd99, 8'd2};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd198, 8'd100, 8'd9};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd209, 8'd108, 8'd20};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd209, 8'd107, 8'd22};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd199, 8'd98, 8'd8};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd191, 8'd94, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd190, 8'd96, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd227, 8'd120, 8'd26};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd250, 8'd152, 8'd61};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd220, 8'd131, 8'd41};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd194, 8'd106, 8'd17};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd176, 8'd89, 8'd9};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd169, 8'd91, 8'd29};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd144, 8'd85, 8'd53};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd138, 8'd96, 8'd84};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd87, 8'd98, 8'd102};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd92, 8'd105, 8'd111};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd140, 8'd159, 8'd166};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd184, 8'd207, 8'd215};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd182, 8'd205, 8'd211};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd173, 8'd197, 8'd199};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd172, 8'd192, 8'd191};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd155, 8'd174, 8'd170};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd178, 8'd185, 8'd154};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd205, 8'd209, 8'd174};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd119, 8'd87, 8'd74};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd111, 8'd68, 8'd52};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd105, 8'd57, 8'd43};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd78, 8'd30, 8'd20};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd49, 8'd2, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd34, 8'd25, 8'd18};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd189, 8'd184, 8'd178};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd192, 8'd210, 8'd210};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd115, 8'd135, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd66, 8'd87, 8'd92};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd85, 8'd108, 8'd114};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd133, 8'd158, 8'd163};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd171, 8'd190, 8'd196};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd195, 8'd213, 8'd217};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd187, 8'd209, 8'd206};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd154, 8'd174, 8'd172};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd169, 8'd188, 8'd186};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd199, 8'd184, 8'd179};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd24, 8'd0, 8'd0};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd58, 8'd21, 8'd13};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd91, 8'd47, 8'd38};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd119, 8'd71, 8'd59};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd126, 8'd77, 8'd63};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd123, 8'd94, 8'd88};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd246, 8'd218, 8'd170};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd238, 8'd215, 8'd174};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd198, 8'd183, 8'd154};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd173, 8'd167, 8'd153};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd185, 8'd190, 8'd186};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd203};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd175, 8'd192, 8'd199};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd181, 8'd202, 8'd207};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd199, 8'd213, 8'd222};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd159, 8'd180, 8'd183};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd116, 8'd142, 8'd139};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd96, 8'd116, 8'd115};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd99, 8'd93, 8'd93};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd116, 8'd74, 8'd58};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd144, 8'd67, 8'd23};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd169, 8'd70, 8'd3};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd189, 8'd95, 8'd0};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd222, 8'd125, 8'd28};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd234, 8'd138, 8'd36};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd237, 8'd139, 8'd38};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd193, 8'd93, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd195, 8'd94, 8'd2};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd203, 8'd99, 8'd14};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd200, 8'd95, 8'd14};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd210, 8'd100, 8'd23};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd195, 8'd93, 8'd11};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd178, 8'd88, 8'd0};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd176, 8'd97, 8'd2};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd193, 8'd122, 8'd18};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd224, 8'd153, 8'd45};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd254, 8'd182, 8'd72};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd87};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd234, 8'd128, 8'd28};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd231, 8'd122, 8'd21};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd234, 8'd121, 8'd17};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd239, 8'd127, 8'd19};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd239, 8'd134, 8'd17};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd235, 8'd141, 8'd17};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd239, 8'd158, 8'd25};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd248, 8'd175, 8'd37};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd246, 8'd172, 8'd23};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd242, 8'd172, 8'd16};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd239, 8'd174, 8'd12};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd238, 8'd179, 8'd25};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd239, 8'd190, 8'd59};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd248, 8'd208, 8'd113};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd172};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd209};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd217};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd174};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd131};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd104};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd241, 8'd210, 8'd104};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd238, 8'd210, 8'd85};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd234, 8'd210, 8'd58};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd234, 8'd212, 8'd41};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd241, 8'd214, 8'd45};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd253, 8'd215, 8'd68};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd96};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd114};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd93};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd74};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd242, 8'd162, 8'd49};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd237, 8'd141, 8'd31};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd25};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd246, 8'd173, 8'd9};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd221, 8'd180, 8'd54};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd174};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd46: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd252, 8'd253, 8'd219};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd247, 8'd202, 8'd99};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd245, 8'd173, 8'd27};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd244, 8'd173, 8'd23};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd0};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd23};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd244, 8'd171, 8'd58};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd246, 8'd187, 8'd87};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd251, 8'd208, 8'd96};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd94};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd252, 8'd218, 8'd84};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd246, 8'd213, 8'd74};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd252, 8'd209, 8'd81};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd93};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd94};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd252, 8'd215, 8'd75};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd237, 8'd206, 8'd56};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd232, 8'd204, 8'd68};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd114};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd157};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd198};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd252, 8'd238, 8'd203};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd249, 8'd238, 8'd216};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd234};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd243};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd234};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd210};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd186};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd243, 8'd188, 8'd95};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd238, 8'd181, 8'd68};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd237, 8'd173, 8'd37};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd246, 8'd173, 8'd18};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd17};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd23};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd252, 8'd159, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd244, 8'd147, 8'd34};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd245, 8'd133, 8'd25};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd243, 8'd128, 8'd22};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd222, 8'd110, 8'd8};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd206, 8'd115, 8'd8};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd249, 8'd184, 8'd68};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd84};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd250, 8'd199, 8'd72};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd247, 8'd188, 8'd62};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd218, 8'd136, 8'd34};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd201, 8'd115, 8'd16};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd188, 8'd95, 8'd2};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd194, 8'd92, 8'd7};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd203, 8'd97, 8'd13};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd205, 8'd96, 8'd11};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd205, 8'd97, 8'd9};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd204, 8'd99, 8'd7};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd201, 8'd93, 8'd5};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd230, 8'd130, 8'd44};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd229, 8'd135, 8'd47};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd205, 8'd110, 8'd18};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd173, 8'd75, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd164, 8'd71, 8'd1};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd136, 8'd61, 8'd19};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd132, 8'd71, 8'd50};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd87, 8'd96, 8'd93};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd97, 8'd109, 8'd109};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd128, 8'd146, 8'd150};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd164, 8'd187, 8'd193};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd179, 8'd204, 8'd211};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd177, 8'd202, 8'd207};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd173, 8'd197, 8'd201};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd172, 8'd193, 8'd196};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd169, 8'd170, 8'd154};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd179, 8'd168, 8'd136};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd201, 8'd174, 8'd121};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd228, 8'd188, 8'd118};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd248, 8'd202, 8'd127};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd253, 8'd214, 8'd145};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd253, 8'd226, 8'd171};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd253, 8'd236, 8'd192};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd147, 8'd120, 8'd111};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd72, 8'd38, 8'd26};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd83, 8'd43, 8'd31};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd62, 8'd22, 8'd14};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd41, 8'd2, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd12, 8'd8, 8'd0};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd121, 8'd121, 8'd113};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd209, 8'd234, 8'd231};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd143, 8'd169, 8'd168};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd71, 8'd101, 8'd103};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd72, 8'd103, 8'd106};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd121, 8'd156, 8'd162};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd131, 8'd168, 8'd176};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd99, 8'd137, 8'd146};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd88, 8'd128, 8'd128};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd95, 8'd134, 8'd133};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd132, 8'd164, 8'd163};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd189, 8'd213, 8'd213};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd179, 8'd203, 8'd205};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd133, 8'd161, 8'd162};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd114, 8'd146, 8'd145};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd101, 8'd135, 8'd134};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd78, 8'd110, 8'd109};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd63, 8'd93, 8'd93};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd68, 8'd96, 8'd97};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd184, 8'd205, 8'd200};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd208, 8'd227, 8'd223};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd124, 8'd106, 8'd102};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd26, 8'd0, 8'd0};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd56, 8'd22, 8'd13};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd71, 8'd33, 8'd20};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd86, 8'd49, 8'd31};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd73, 8'd38, 8'd18};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd166, 8'd145, 8'd128};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd210};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd254, 8'd234, 8'd181};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd249, 8'd220, 8'd152};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd242, 8'd207, 8'd126};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd238, 8'd198, 8'd111};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd217, 8'd165, 8'd89};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd199, 8'd163, 8'd101};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd164, 8'd150, 8'd113};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd160, 8'd166, 8'd154};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd187, 8'd207, 8'd208};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd188, 8'd211, 8'd217};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd178, 8'd198, 8'd199};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd191, 8'd207, 8'd204};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd185, 8'd195, 8'd207};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd144, 8'd162, 8'd166};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd108, 8'd130, 8'd128};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd96, 8'd110, 8'd110};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd100, 8'd86, 8'd85};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd114, 8'd58, 8'd41};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd146, 8'd54, 8'd7};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd184, 8'd67, 8'd0};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd198, 8'd99, 8'd6};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd227, 8'd128, 8'd35};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd236, 8'd135, 8'd43};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd210, 8'd106, 8'd17};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd197, 8'd89, 8'd1};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd208, 8'd97, 8'd15};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd202, 8'd89, 8'd9};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd200, 8'd87, 8'd7};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd185, 8'd80, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd185, 8'd90, 8'd0};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd193, 8'd115, 8'd15};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd216, 8'd154, 8'd41};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd242, 8'd192, 8'd67};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd78};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd69};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd249, 8'd198, 8'd57};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd235, 8'd135, 8'd23};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd227, 8'd123, 8'd10};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd227, 8'd117, 8'd4};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd240, 8'd129, 8'd13};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd248, 8'd144, 8'd21};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd247, 8'd156, 8'd26};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd28};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd244, 8'd175, 8'd35};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd242, 8'd167, 8'd22};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd236, 8'd169, 8'd36};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd231, 8'd178, 8'd62};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd237, 8'd200, 8'd109};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd251, 8'd226, 8'd159};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd203};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd227};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd236};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd224};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd208};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd247, 8'd234, 8'd181};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd236, 8'd220, 8'd145};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd231, 8'd208, 8'd114};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd235, 8'd203, 8'd90};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd245, 8'd206, 8'd79};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd254, 8'd210, 8'd77};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd249, 8'd205, 8'd82};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd253, 8'd214, 8'd83};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd82};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd253, 8'd222, 8'd79};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd245, 8'd216, 8'd78};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd246, 8'd210, 8'd88};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd252, 8'd211, 8'd106};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd123};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd71};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd239, 8'd175, 8'd43};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd239, 8'd156, 8'd34};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd247, 8'd151, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd14};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd240, 8'd171, 8'd6};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd227, 8'd191, 8'd81};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd214};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd47: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd225};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd248, 8'd210, 8'd109};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd36};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd244, 8'd178, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd3};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd248, 8'd163, 8'd10};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd240, 8'd148, 8'd25};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd250, 8'd159, 8'd54};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd85};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd110};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd118};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd242, 8'd220, 8'd118};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd71};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd251, 8'd215, 8'd92};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd109};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd102};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd252, 8'd214, 8'd81};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd69};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd207, 8'd77};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd241, 8'd205, 8'd93};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd235, 8'd206, 8'd102};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd245, 8'd212, 8'd115};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd138};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd164};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd190};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd217};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd243};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd247, 8'd255, 8'd251};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd190};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd253, 8'd214, 8'd139};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd235, 8'd185, 8'd70};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd235, 8'd174, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd252, 8'd174, 8'd12};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd18};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd24};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd249, 8'd137, 8'd25};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd251, 8'd146, 8'd31};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd236, 8'd128, 8'd17};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd210, 8'd108, 8'd0};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd202, 8'd120, 8'd8};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd244, 8'd190, 8'd68};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd245, 8'd206, 8'd75};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd76};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd90};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd106};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd247, 8'd165, 8'd65};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd202, 8'd111, 8'd18};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd184, 8'd82, 8'd0};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd186, 8'd77, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd192, 8'd80, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd198, 8'd86, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd203, 8'd92, 8'd3};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd201, 8'd95, 8'd7};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd206, 8'd106, 8'd18};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd225, 8'd130, 8'd36};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd225, 8'd127, 8'd28};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd185, 8'd83, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd168, 8'd69, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd132, 8'd49, 8'd0};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd124, 8'd53, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd91, 8'd101, 8'd93};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd106, 8'd118, 8'd114};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd115, 8'd133, 8'd133};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd141, 8'd165, 8'd169};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd178, 8'd205, 8'd212};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd183, 8'd210, 8'd219};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd175, 8'd200, 8'd207};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd185, 8'd210, 8'd217};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd197, 8'd189, 8'd187};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd180, 8'd156, 8'd132};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd176, 8'd127, 8'd68};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd194, 8'd128, 8'd34};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd216, 8'd146, 8'd35};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd226, 8'd165, 8'd58};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd228, 8'd188, 8'd92};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd233, 8'd206, 8'd119};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd194, 8'd171, 8'd163};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd60, 8'd30, 8'd19};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd64, 8'd32, 8'd21};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd54, 8'd20, 8'd11};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd53, 8'd20, 8'd15};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd22, 8'd19, 8'd10};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd68, 8'd69, 8'd61};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd194, 8'd199, 8'd195};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd225, 8'd230, 8'd224};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd129, 8'd160, 8'd155};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd92, 8'd122, 8'd120};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd76, 8'd110, 8'd109};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd99, 8'd137, 8'd138};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd120, 8'd159, 8'd164};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd111, 8'd154, 8'd161};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd102, 8'd149, 8'd157};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd110, 8'd157, 8'd167};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd104, 8'd159, 8'd156};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd85, 8'd135, 8'd132};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd71, 8'd113, 8'd111};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd93, 8'd125, 8'd122};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd156, 8'd178, 8'd175};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd223, 8'd235, 8'd231};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd128, 8'd156, 8'd160};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd93, 8'd124, 8'd127};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd94, 8'd129, 8'd131};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd116, 8'd156, 8'd156};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd112, 8'd154, 8'd153};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd104, 8'd144, 8'd144};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd102, 8'd140, 8'd141};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd95, 8'd130, 8'd132};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd66, 8'd95, 8'd90};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd116, 8'd141, 8'd137};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd181, 8'd201, 8'd199};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd223, 8'd215, 8'd212};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd57, 8'd39, 8'd35};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd34, 8'd7, 8'd0};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd45, 8'd13, 8'd2};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd65, 8'd33, 8'd18};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd84, 8'd56, 8'd35};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd69, 8'd43, 8'd20};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd200, 8'd182, 8'd160};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd251, 8'd229, 8'd179};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd245, 8'd210, 8'd129};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd233, 8'd186, 8'd78};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd221, 8'd166, 8'd37};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd214, 8'd155, 8'd15};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd191, 8'd127, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd154, 8'd108, 8'd33};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd154, 8'd141, 8'd99};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd177, 8'd190, 8'd180};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd172, 8'd203, 8'd208};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd174, 8'd204, 8'd212};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd192, 8'd214, 8'd212};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd197, 8'd210, 8'd201};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd163, 8'd169, 8'd183};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd132, 8'd145, 8'd153};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd104, 8'd122, 8'd122};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd97, 8'd107, 8'd108};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd99, 8'd79, 8'd78};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd113, 8'd52, 8'd34};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd156, 8'd54, 8'd6};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd203, 8'd75, 8'd4};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd199, 8'd99, 8'd11};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd217, 8'd116, 8'd28};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd221, 8'd117, 8'd32};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd181, 8'd72, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd203, 8'd90, 8'd10};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd201, 8'd86, 8'd6};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd182, 8'd65, 8'd0};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd198, 8'd78, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd197, 8'd96, 8'd4};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd222, 8'd133, 8'd33};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd251, 8'd181, 8'd69};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd86};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd79};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd247, 8'd217, 8'd59};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd238, 8'd206, 8'd43};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd234, 8'd199, 8'd33};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd233, 8'd134, 8'd14};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd229, 8'd124, 8'd6};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd234, 8'd123, 8'd5};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd137, 8'd17};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd24};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd250, 8'd156, 8'd24};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd241, 8'd159, 8'd21};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd23};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd244, 8'd166, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd251, 8'd185, 8'd75};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd145};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd205};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd237};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd251, 8'd251, 8'd241};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd246, 8'd251, 8'd229};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd244, 8'd251, 8'd218};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd246, 8'd221, 8'd154};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd244, 8'd217, 8'd136};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd241, 8'd214, 8'd109};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd244, 8'd215, 8'd89};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd249, 8'd218, 8'd76};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd253, 8'd218, 8'd74};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd251, 8'd216, 8'd74};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd74};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd83};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd86};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd254, 8'd211, 8'd96};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd253, 8'd216, 8'd110};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd122};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd128};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd126};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd122};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd243, 8'd185, 8'd39};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd229, 8'd165, 8'd16};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd27};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd252, 8'd160, 8'd0};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd244, 8'd179, 8'd15};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd117};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd48: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd250, 8'd205, 8'd90};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd236, 8'd171, 8'd0};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd249, 8'd171, 8'd23};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd17};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd6};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd233, 8'd149, 8'd15};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd238, 8'd157, 8'd65};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd123};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd142};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd253, 8'd222, 8'd131};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd246, 8'd225, 8'd118};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd254, 8'd226, 8'd117};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd105};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd88};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd87};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd98};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd251, 8'd218, 8'd105};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd242, 8'd214, 8'd104};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd71};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd252, 8'd211, 8'd67};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd245, 8'd208, 8'd65};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd241, 8'd207, 8'd73};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd241, 8'd210, 8'd93};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd246, 8'd218, 8'd121};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd151};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd170};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd234};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd223};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd192};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd237, 8'd230, 8'd140};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd218, 8'd197, 8'd80};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd213, 8'd171, 8'd35};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd222, 8'd161, 8'd11};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd234, 8'd159, 8'd5};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd249, 8'd157, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd236, 8'd143, 8'd14};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd229, 8'd132, 8'd2};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd222, 8'd125, 8'd0};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd248, 8'd160, 8'd26};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd56};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd254, 8'd188, 8'd50};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd67};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd87};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd247, 8'd219, 8'd86};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd246, 8'd215, 8'd90};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd242, 8'd201, 8'd85};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd222, 8'd163, 8'd61};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd196, 8'd112, 8'd26};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd182, 8'd74, 8'd2};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd182, 8'd60, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd187, 8'd67, 8'd4};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd197, 8'd79, 8'd17};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd206, 8'd91, 8'd26};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd204, 8'd94, 8'd17};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd188, 8'd83, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd170, 8'd66, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd156, 8'd51, 8'd3};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd152, 8'd44, 8'd18};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd112, 8'd69, 8'd86};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd102, 8'd99, 8'd108};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd95, 8'd127, 8'd126};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd111, 8'd147, 8'd135};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd161, 8'd174, 8'd157};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd201, 8'd203, 8'd190};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd194, 8'd215, 8'd210};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd164, 8'd210, 8'd210};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd169, 8'd208, 8'd190};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd180, 8'd193, 8'd176};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd163, 8'd136, 8'd107};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd156, 8'd94, 8'd37};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd194, 8'd111, 8'd15};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd205, 8'd117, 8'd0};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd242, 8'd156, 8'd17};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd29};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd247, 8'd192, 8'd91};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd125};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd177};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd218};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd13, 8'd18, 8'd14};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd34, 8'd40, 8'd36};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd59, 8'd68, 8'd63};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd63, 8'd74, 8'd68};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd79, 8'd105, 8'd104};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd75, 8'd101, 8'd100};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd100, 8'd124, 8'd124};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd208, 8'd234, 8'd233};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd195, 8'd224, 8'd222};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd160, 8'd192, 8'd189};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd105, 8'd141, 8'd137};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd74, 8'd113, 8'd108};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd69, 8'd118, 8'd115};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd96, 8'd145, 8'd142};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd116, 8'd165, 8'd162};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd113, 8'd162, 8'd159};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd100, 8'd149, 8'd146};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd91, 8'd141, 8'd138};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd86, 8'd136, 8'd133};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd80, 8'd130, 8'd127};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd71, 8'd118, 8'd108};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd82, 8'd125, 8'd116};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd86, 8'd126, 8'd118};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd81, 8'd113, 8'd108};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd82, 8'd108, 8'd105};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd120, 8'd138, 8'd138};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd192, 8'd206, 8'd207};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd156, 8'd174, 8'd176};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd66, 8'd85, 8'd89};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd72, 8'd107, 8'd113};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd83, 8'd120, 8'd126};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd99, 8'd138, 8'd143};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd105, 8'd149, 8'd152};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd103, 8'd151, 8'd153};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd100, 8'd151, 8'd152};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd99, 8'd153, 8'd153};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd101, 8'd157, 8'd156};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd108, 8'd154, 8'd152};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd83, 8'd127, 8'd126};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd72, 8'd111, 8'd110};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd95, 8'd126, 8'd128};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd148, 8'd172, 8'd174};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd209, 8'd227, 8'd231};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd229, 8'd232, 8'd237};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd128, 8'd132, 8'd135};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd69, 8'd74, 8'd77};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd55, 8'd56, 8'd58};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd42, 8'd36, 8'd40};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd45, 8'd28, 8'd34};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd63, 8'd33, 8'd41};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd87, 8'd49, 8'd60};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd248, 8'd207, 8'd153};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd121};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd249, 8'd194, 8'd75};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd243, 8'd179, 8'd45};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd233, 8'd160, 8'd29};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd194, 8'd115, 8'd0};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd182, 8'd100, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd187, 8'd82, 8'd14};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd175, 8'd122, 8'd72};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd181, 8'd184, 8'd163};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd177, 8'd202, 8'd207};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd194, 8'd209, 8'd228};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd192, 8'd199, 8'd217};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd189, 8'd212, 8'd220};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd164, 8'd208, 8'd207};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd130, 8'd146, 8'd169};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd102, 8'd128, 8'd141};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd96, 8'd122, 8'd123};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd94};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd104, 8'd66, 8'd43};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd128, 8'd49, 8'd10};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd167, 8'd62, 8'd7};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd186, 8'd71, 8'd6};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd196, 8'd97, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd187, 8'd78, 8'd13};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd186, 8'd62, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd190, 8'd61, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd189, 8'd67, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd186, 8'd85, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd201, 8'd123, 8'd22};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd222, 8'd160, 8'd51};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd84};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd78};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd80};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd253, 8'd219, 8'd70};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd237, 8'd197, 8'd50};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd242, 8'd193, 8'd52};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd62};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd253, 8'd191, 8'd58};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd236, 8'd127, 8'd24};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd233, 8'd132, 8'd14};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd230, 8'd140, 8'd2};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd225, 8'd150, 8'd0};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd221, 8'd160, 8'd7};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd224, 8'd173, 8'd32};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd230, 8'd186, 8'd63};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd235, 8'd193, 8'd81};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd251, 8'd239, 8'd189};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd197};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd202};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd196};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd171};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd131};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd248, 8'd212, 8'd89};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd242, 8'd205, 8'd62};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd223, 8'd214, 8'd77};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd233, 8'd217, 8'd82};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd245, 8'd221, 8'd87};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd91};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd92};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd92};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd92};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd246, 8'd209, 8'd92};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd250, 8'd202, 8'd76};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd254, 8'd218, 8'd106};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd244, 8'd223, 8'd134};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd230, 8'd218, 8'd144};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd237, 8'd218, 8'd149};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd136};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd93};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd244, 8'd163, 8'd48};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd15};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd245, 8'd160, 8'd18};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd240, 8'd169, 8'd19};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd248, 8'd174, 8'd15};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd253, 8'd172, 8'd20};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd248, 8'd182, 8'd70};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd245, 8'd217, 8'd169};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd49: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd251, 8'd212, 8'd117};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd239, 8'd183, 8'd34};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd253, 8'd178, 8'd11};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd18};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd27};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd250, 8'd159, 8'd29};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd237, 8'd152, 8'd35};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd234, 8'd163, 8'd57};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd251, 8'd196, 8'd105};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd146};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd251, 8'd234, 8'd142};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd239, 8'd219, 8'd124};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd114};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd119};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd116};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd213, 8'd99};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd249, 8'd208, 8'd90};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd95};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd98};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd94};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd254, 8'd217, 8'd87};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd249, 8'd214, 8'd84};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd245, 8'd213, 8'd90};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd244, 8'd212, 8'd101};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd114};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd243, 8'd212, 8'd122};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd247, 8'd223, 8'd127};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd251, 8'd229, 8'd146};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd175};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd195};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd187};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd149};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd237, 8'd186, 8'd94};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd218, 8'd160, 8'd52};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd228, 8'd150, 8'd26};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd223, 8'd143, 8'd20};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd217, 8'd133, 8'd8};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd212, 8'd129, 8'd1};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd235, 8'd158, 8'd26};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd53};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd243, 8'd190, 8'd48};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd232, 8'd186, 8'd41};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd250, 8'd215, 8'd69};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd80};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd90};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd91};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd88};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd251, 8'd187, 8'd81};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd239, 8'd156, 8'd62};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd222, 8'd128, 8'd40};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd178, 8'd75, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd174, 8'd71, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd175, 8'd72, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd182, 8'd81, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd188, 8'd90, 8'd3};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd180, 8'd80, 8'd5};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd157, 8'd55, 8'd6};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd139, 8'd33, 8'd7};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd108, 8'd57, 8'd62};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd106, 8'd94, 8'd96};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd96, 8'd124, 8'd125};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd100, 8'd136, 8'd132};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd141, 8'd160, 8'd154};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd191, 8'd196, 8'd190};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd197, 8'd213, 8'd212};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd171, 8'd206, 8'd208};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd179, 8'd211, 8'd206};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd186, 8'd205, 8'd201};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd172, 8'd158, 8'd145};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd167, 8'd113, 8'd77};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd179, 8'd88, 8'd18};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd200, 8'd98, 8'd0};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd222, 8'd132, 8'd12};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd234, 8'd159, 8'd32};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd246, 8'd176, 8'd54};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd241, 8'd181, 8'd71};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd235, 8'd194, 8'd106};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd238, 8'd213, 8'd149};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd248, 8'd233, 8'd192};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd77};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd78, 8'd92, 8'd92};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd100, 8'd116, 8'd116};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd101, 8'd119, 8'd119};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd80, 8'd108, 8'd109};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd82, 8'd110, 8'd111};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd82, 8'd112, 8'd112};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd117, 8'd147, 8'd147};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd98, 8'd130, 8'd129};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd83, 8'd119, 8'd117};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd97, 8'd136, 8'd133};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd113, 8'd154, 8'd150};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd133, 8'd179, 8'd177};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd121, 8'd167, 8'd165};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd110, 8'd154, 8'd153};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd104, 8'd148, 8'd147};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd102, 8'd144, 8'd143};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd94, 8'd134, 8'd134};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd81, 8'd121, 8'd121};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd73, 8'd111, 8'd112};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd66, 8'd103, 8'd96};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd36, 8'd71, 8'd65};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd30, 8'd61, 8'd56};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd47, 8'd73, 8'd70};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd45, 8'd67, 8'd65};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd50, 8'd66, 8'd66};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd114, 8'd128, 8'd129};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd199, 8'd210, 8'd212};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd224, 8'd232, 8'd235};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd156, 8'd167, 8'd171};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd101, 8'd116, 8'd119};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd102};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd69, 8'd100, 8'd105};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd75, 8'd106, 8'd111};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd79, 8'd114, 8'd118};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd83, 8'd121, 8'd124};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd87, 8'd128, 8'd130};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd92, 8'd136, 8'd137};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd97, 8'd145, 8'd145};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd102, 8'd150, 8'd150};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd105, 8'd149, 8'd150};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd116, 8'd157, 8'd159};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd108, 8'd146, 8'd147};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd97, 8'd131, 8'd133};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd92, 8'd121, 8'd125};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd91, 8'd116, 8'd120};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd121, 8'd142, 8'd147};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd173, 8'd192, 8'd198};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd159, 8'd180, 8'd181};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd99, 8'd123, 8'd123};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd81, 8'd105, 8'd105};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd86, 8'd108, 8'd106};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd73, 8'd87, 8'd87};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd74, 8'd78, 8'd81};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd69, 8'd63, 8'd67};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd100, 8'd87, 8'd94};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd240, 8'd189, 8'd126};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd236, 8'd181, 8'd101};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd246, 8'd183, 8'd80};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd249, 8'd177, 8'd56};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd245, 8'd163, 8'd38};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd227, 8'd137, 8'd25};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd200, 8'd103, 8'd9};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd191, 8'd90, 8'd10};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd179, 8'd81, 8'd20};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd154, 8'd102, 8'd62};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd168, 8'd170, 8'd156};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd183, 8'd208, 8'd215};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd188, 8'd204, 8'd219};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd198, 8'd202, 8'd213};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd195, 8'd209, 8'd209};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd153, 8'd185, 8'd174};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd117, 8'd138, 8'd157};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd99, 8'd123, 8'd135};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd94, 8'd112, 8'd112};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd100, 8'd90, 8'd78};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd105, 8'd55, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd131, 8'd46, 8'd5};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd167, 8'd64, 8'd5};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd182, 8'd75, 8'd3};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd197, 8'd106, 8'd27};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd172, 8'd76, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd162, 8'd61, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd189, 8'd89, 8'd4};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd230, 8'd137, 8'd44};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd254, 8'd175, 8'd74};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd90};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd96};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd254, 8'd217, 8'd84};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd84};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd82};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd248, 8'd212, 8'd64};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd241, 8'd199, 8'd53};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd250, 8'd199, 8'd56};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd250, 8'd191, 8'd53};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd235, 8'd171, 8'd37};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd228, 8'd142, 8'd0};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd230, 8'd151, 8'd0};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd231, 8'd158, 8'd3};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd224, 8'd162, 8'd19};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd222, 8'd167, 8'd50};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd233, 8'd186, 8'd98};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd155};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd196};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd154};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd151};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd245, 8'd219, 8'd142};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd240, 8'd208, 8'd131};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd239, 8'd205, 8'd118};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd245, 8'd207, 8'd106};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd254, 8'd215, 8'd98};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd93};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd250, 8'd223, 8'd90};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd251, 8'd221, 8'd89};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd90};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd92};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd254, 8'd212, 8'd94};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd102};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd110};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd117};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd115};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd245, 8'd213, 8'd112};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd245, 8'd220, 8'd130};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd157};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd144};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd237, 8'd188, 8'd93};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd233, 8'd165, 8'd54};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd46};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd17};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd17};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd10};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd244, 8'd170, 8'd13};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd247, 8'd179, 8'd44};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd251, 8'd204, 8'd112};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd198};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd50: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd252, 8'd227, 8'd163};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd245, 8'd204, 8'd98};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd10};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd20};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd32};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd249, 8'd161, 8'd12};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd235, 8'd159, 8'd14};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd242, 8'd174, 8'd63};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd118};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd247, 8'd225, 8'd140};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd249, 8'd228, 8'd145};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd249, 8'd228, 8'd147};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd246, 8'd224, 8'd139};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd247, 8'd221, 8'd128};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd253, 8'd219, 8'd112};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd98};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd86};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd119};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd114};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd105};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd97};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd252, 8'd217, 8'd91};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd247, 8'd212, 8'd86};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd242, 8'd206, 8'd86};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd238, 8'd201, 8'd84};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd74};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd246, 8'd199, 8'd81};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd234, 8'd194, 8'd99};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd236, 8'd202, 8'd130};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd155};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd162};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd148};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd131};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd250, 8'd187, 8'd73};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd247, 8'd180, 8'd65};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd228, 8'd155, 8'd40};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd215, 8'd143, 8'd22};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd221, 8'd153, 8'd26};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd241, 8'd183, 8'd47};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd248, 8'd203, 8'd58};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd223, 8'd186, 8'd36};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd238, 8'd193, 8'd38};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd58};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd75};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd80};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd85};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd92};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd94};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd91};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd85};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd232, 8'd151, 8'd59};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd194, 8'd110, 8'd20};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd171, 8'd86, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd167, 8'd80, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd165, 8'd73, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd154, 8'd57, 8'd6};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd144, 8'd40, 8'd13};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd111, 8'd45, 8'd29};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd111, 8'd86, 8'd79};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd98, 8'd118, 8'd119};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd88, 8'd125, 8'd133};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd118, 8'd145, 8'd152};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd173, 8'd184, 8'd188};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd211};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd186, 8'd205, 8'd211};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd179, 8'd204, 8'd211};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd181, 8'd208, 8'd215};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd178, 8'd188, 8'd189};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd182, 8'd140, 8'd126};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd170, 8'd71, 8'd32};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd203, 8'd80, 8'd13};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd205, 8'd105, 8'd11};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd214, 8'd144, 8'd33};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd250, 8'd164, 8'd19};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd248, 8'd167, 8'd32};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd241, 8'd174, 8'd59};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd236, 8'd183, 8'd87};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd236, 8'd193, 8'd115};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd240, 8'd200, 8'd138};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd245, 8'd205, 8'd153};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd248, 8'd208, 8'd157};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd105, 8'd124, 8'd128};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd95, 8'd118, 8'd124};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd83, 8'd110, 8'd117};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd62, 8'd91, 8'd99};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd78, 8'd112, 8'd114};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd102, 8'd136, 8'd138};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd111, 8'd146, 8'd148};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd117, 8'd155, 8'd156};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd135, 8'd173, 8'd174};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd132, 8'd172, 8'd172};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd140, 8'd180, 8'd180};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd137, 8'd177, 8'd177};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd108, 8'd150, 8'd148};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd109, 8'd149, 8'd148};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd111, 8'd150, 8'd149};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd108, 8'd142, 8'd143};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd93, 8'd123, 8'd125};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd86, 8'd111, 8'd115};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd105, 8'd129, 8'd133};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd136, 8'd157, 8'd162};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd167, 8'd187, 8'd185};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd176, 8'd196, 8'd194};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd203, 8'd222, 8'd220};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd205, 8'd219, 8'd219};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd210, 8'd222, 8'd222};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd187, 8'd192, 8'd196};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd124, 8'd134, 8'd136};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd99, 8'd113, 8'd116};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd110, 8'd124, 8'd127};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd126, 8'd146, 8'd153};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd108, 8'd131, 8'd137};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd87, 8'd112, 8'd117};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd72, 8'd100, 8'd104};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd73, 8'd102, 8'd106};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd83, 8'd117, 8'd119};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd98, 8'd133, 8'd135};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd108, 8'd143, 8'd145};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd113, 8'd151, 8'd154};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd110, 8'd148, 8'd151};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd165, 8'd168};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd129, 8'd167, 8'd170};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd105, 8'd143, 8'd146};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd105, 8'd143, 8'd146};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd112, 8'd150, 8'd153};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd96, 8'd131, 8'd135};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd82, 8'd128, 8'd126};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd69, 8'd115, 8'd112};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd83, 8'd128, 8'd125};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd84, 8'd126, 8'd122};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd80, 8'd116, 8'd114};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd91, 8'd120, 8'd118};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd78, 8'd100, 8'd98};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd121, 8'd139, 8'd139};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd197, 8'd163, 8'd136};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd194, 8'd150, 8'd111};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd193, 8'd142, 8'd89};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd196, 8'd138, 8'd74};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd196, 8'd136, 8'd64};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd228, 8'd159, 8'd64};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd233, 8'd160, 8'd55};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd239, 8'd158, 8'd41};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd40};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd239, 8'd139, 8'd27};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd206, 8'd97, 8'd6};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd190, 8'd75, 8'd8};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd182, 8'd65, 8'd12};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd174, 8'd75, 8'd18};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd136, 8'd82, 8'd44};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd151, 8'd147, 8'd136};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd188, 8'd208, 8'd215};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd183, 8'd201, 8'd213};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd201, 8'd209, 8'd212};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd188, 8'd199, 8'd193};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd132, 8'd154, 8'd141};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd107, 8'd131, 8'd143};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd102, 8'd121, 8'd127};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd103, 8'd105, 8'd102};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd104, 8'd75, 8'd61};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd113, 8'd46, 8'd19};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd143, 8'd52, 8'd7};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd173, 8'd78, 8'd12};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd183, 8'd92, 8'd11};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd159, 8'd80, 8'd0};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd190, 8'd116, 8'd17};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd236, 8'd169, 8'd65};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd102};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd107};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd92};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd248, 8'd208, 8'd86};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd253, 8'd213, 8'd91};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd254, 8'd214, 8'd83};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd91};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd251, 8'd212, 8'd73};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd237, 8'd196, 8'd52};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd245, 8'd199, 8'd54};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd60};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd244, 8'd180, 8'd44};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd224, 8'd156, 8'd23};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd226, 8'd151, 8'd24};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd229, 8'd157, 8'd36};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd238, 8'd173, 8'd57};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd193, 8'd86};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd114};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd128};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd245, 8'd213, 8'd128};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd233, 8'd207, 8'd123};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd251, 8'd220, 8'd103};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd247, 8'd217, 8'd97};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd241, 8'd209, 8'd90};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd238, 8'd203, 8'd85};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd240, 8'd203, 8'd88};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd245, 8'd208, 8'd94};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd254, 8'd214, 8'd103};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd110};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd92};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd88};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd254, 8'd209, 8'd90};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd101};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd116};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd129};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd254, 8'd226, 8'd129};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd245, 8'd222, 8'd128};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd252, 8'd228, 8'd140};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd145};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd144};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd127};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd246, 8'd193, 8'd89};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd230, 8'd167, 8'd51};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd234, 8'd161, 8'd33};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd246, 8'd168, 8'd32};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd20};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd9};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd1};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd244, 8'd170, 8'd21};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd239, 8'd195, 8'd86};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd253, 8'd233, 8'd174};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd51: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd252, 8'd242, 8'd207};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd250, 8'd224, 8'd165};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd245, 8'd181, 8'd32};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd248, 8'd175, 8'd34};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd29};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd19};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd9};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd15};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd243, 8'd164, 8'd37};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd239, 8'd161, 8'd60};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd240, 8'd191, 8'd98};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd129};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd156};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd249, 8'd229, 8'd156};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd240, 8'd223, 8'd145};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd246, 8'd225, 8'd134};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd118};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd250, 8'd217, 8'd102};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd244, 8'd209, 8'd117};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd114};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd107};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd252, 8'd217, 8'd99};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd94};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd91};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd213, 8'd89};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd252, 8'd210, 8'd89};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd95};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd88};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd247, 8'd204, 8'd74};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd233, 8'd199, 8'd65};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd226, 8'd196, 8'd62};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd226, 8'd197, 8'd69};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd233, 8'd201, 8'd82};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd240, 8'd204, 8'd92};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd98};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd89};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd241, 8'd168, 8'd65};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd234, 8'd160, 8'd51};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd223, 8'd152, 8'd34};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd233, 8'd170, 8'd41};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd70};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd246, 8'd202, 8'd53};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd241, 8'd185, 8'd36};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd238, 8'd188, 8'd39};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd242, 8'd202, 8'd53};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd249, 8'd219, 8'd73};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd246, 8'd223, 8'd81};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd240, 8'd221, 8'd83};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd245, 8'd225, 8'd92};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd104};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd107};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd98};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd240, 8'd178, 8'd77};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd215, 8'd147, 8'd48};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd193, 8'd119, 8'd22};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd174, 8'd92, 8'd10};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd158, 8'd67, 8'd12};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd150, 8'd53, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd123, 8'd45, 8'd9};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd117, 8'd76, 8'd58};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd101, 8'd106, 8'd109};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd88, 8'd121, 8'd136};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd106, 8'd138, 8'd153};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd148, 8'd166, 8'd176};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd185, 8'd194, 8'd201};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd199, 8'd206, 8'd214};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd175, 8'd193, 8'd203};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd163, 8'd198, 8'd204};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd176, 8'd204, 8'd205};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd181, 8'd151, 8'd143};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd177, 8'd73, 8'd48};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd209, 8'd72, 8'd20};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd199, 8'd93, 8'd9};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd193, 8'd128, 8'd24};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd253, 8'd162, 8'd11};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd21};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd250, 8'd169, 8'd38};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd239, 8'd168, 8'd52};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd229, 8'd164, 8'd64};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd219, 8'd159, 8'd73};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd213, 8'd155, 8'd81};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd212, 8'd155, 8'd84};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd221, 8'd186, 8'd144};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd225, 8'd195, 8'd157};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd235, 8'd212, 8'd180};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd188, 8'd212, 8'd214};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd85, 8'd114, 8'd120};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd60, 8'd92, 8'd103};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd63, 8'd101, 8'd114};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd66, 8'd105, 8'd120};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd77, 8'd114, 8'd120};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd133, 8'd172, 8'd177};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd148, 8'd189, 8'd193};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd124, 8'd168, 8'd171};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd125, 8'd169, 8'd172};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd115, 8'd159, 8'd162};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd109, 8'd150, 8'd154};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd107, 8'd146, 8'd151};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd109, 8'd144, 8'd140};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd88, 8'd120, 8'd117};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd81, 8'd110, 8'd108};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd112, 8'd136, 8'd136};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd166, 8'd184, 8'd186};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd226};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd217, 8'd230, 8'd236};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd218, 8'd231, 8'd237};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd218, 8'd233, 8'd238};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd213, 8'd228, 8'd233};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd191, 8'd209, 8'd213};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd152, 8'd171, 8'd175};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd105, 8'd126, 8'd129};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd73, 8'd94, 8'd97};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd79, 8'd108, 8'd114};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd102, 8'd133, 8'd138};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd99, 8'd132, 8'd137};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd108, 8'd145, 8'd151};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd144, 8'd185, 8'd189};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd141, 8'd186, 8'd191};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd113, 8'd162, 8'd166};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd114, 8'd163, 8'd167};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd121, 8'd175, 8'd175};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd115, 8'd167, 8'd165};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd102, 8'd154, 8'd152};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd42, 8'd91, 8'd88};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd44, 8'd90, 8'd88};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd72, 8'd112, 8'd111};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd79, 8'd115, 8'd113};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd128, 8'd162, 8'd161};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd204, 8'd164, 8'd139};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd197, 8'd153, 8'd126};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd188, 8'd135, 8'd103};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd181, 8'd119, 8'd78};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd178, 8'd111, 8'd59};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd181, 8'd110, 8'd46};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd188, 8'd114, 8'd41};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd194, 8'd118, 8'd40};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd208, 8'd131, 8'd27};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd224, 8'd142, 8'd32};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd227, 8'd140, 8'd24};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd245, 8'd150, 8'd34};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd227, 8'd125, 8'd17};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd186, 8'd78, 8'd0};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd181, 8'd68, 8'd0};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd175, 8'd62, 8'd6};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd179, 8'd67, 8'd1};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd145, 8'd74, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd142, 8'd123, 8'd108};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd181, 8'd194, 8'd200};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd179, 8'd201, 8'd212};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd190, 8'd209, 8'd213};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd157, 8'd176, 8'd174};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd111, 8'd132, 8'd127};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd107, 8'd122, 8'd127};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd111, 8'd120, 8'd117};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd114, 8'd100, 8'd89};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd114, 8'd66, 8'd46};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd130, 8'd47, 8'd15};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd161, 8'd65, 8'd14};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd186, 8'd98, 8'd26};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd192, 8'd116, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd226, 8'd164, 8'd55};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd236, 8'd183, 8'd69};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd244, 8'd208, 8'd88};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd242, 8'd218, 8'd92};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd232, 8'd215, 8'd83};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd231, 8'd212, 8'd81};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd246, 8'd222, 8'd90};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd102};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd83};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd82};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd240, 8'd194, 8'd57};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd231, 8'd184, 8'd44};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd250, 8'd197, 8'd55};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd57};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd236, 8'd168, 8'd35};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd226, 8'd151, 8'd23};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd232, 8'd150, 8'd76};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd247, 8'd169, 8'd97};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd188, 8'd116};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd252, 8'd191, 8'd111};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd231, 8'd180, 8'd88};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd215, 8'd178, 8'd63};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd218, 8'd190, 8'd54};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd227, 8'd205, 8'd57};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd248, 8'd201, 8'd85};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd206, 8'd83};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd82};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd82};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd88};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd96};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd252, 8'd214, 8'd103};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd108};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd252, 8'd207, 8'd82};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd253, 8'd208, 8'd89};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd253, 8'd213, 8'd102};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd253, 8'd218, 8'd116};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd129};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd249, 8'd228, 8'd137};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd245, 8'd231, 8'd142};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd242, 8'd232, 8'd143};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd245, 8'd227, 8'd155};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd155};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd122};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd239, 8'd176, 8'd70};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd231, 8'd160, 8'd36};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd248, 8'd170, 8'd34};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd251, 8'd175, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd240, 8'd166, 8'd17};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd251, 8'd177, 8'd18};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd4};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd6};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd249, 8'd184, 8'd56};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd244, 8'd221, 8'd145};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd249, 8'd254, 8'd224};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd52: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd254, 8'd239, 8'd216};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd237, 8'd186, 8'd94};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd244, 8'd185, 8'd65};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd254, 8'd185, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd14};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd14};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd23};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd248, 8'd162, 8'd27};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd244, 8'd164, 8'd27};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd247, 8'd163, 8'd49};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd243, 8'd170, 8'd67};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd249, 8'd195, 8'd107};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd151};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd167};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd245, 8'd232, 8'd154};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd227, 8'd142};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd249, 8'd234, 8'd141};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd243, 8'd216, 8'd111};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd244, 8'd216, 8'd109};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd245, 8'd215, 8'd105};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd247, 8'd214, 8'd101};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd251, 8'd215, 8'd101};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd103};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd106};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd108};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd251, 8'd207, 8'd98};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd100};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd96};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd82};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd243, 8'd205, 8'd60};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd229, 8'd186, 8'd47};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd225, 8'd176, 8'd47};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd225, 8'd173, 8'd51};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd228, 8'd158, 8'd63};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd231, 8'd156, 8'd63};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd235, 8'd152, 8'd60};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd250, 8'd163, 8'd68};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd234, 8'd149, 8'd43};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd226, 8'd150, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd61};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd63};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd64};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd243, 8'd185, 8'd49};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd231, 8'd183, 8'd47};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd241, 8'd205, 8'd69};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd93};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd104};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd244, 8'd229, 8'd100};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd237, 8'd224, 8'd96};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd246, 8'd213, 8'd82};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd92};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd246, 8'd202, 8'd95};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd233, 8'd180, 8'd78};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd208, 8'd146, 8'd47};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd180, 8'd108, 8'd23};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd159, 8'd77, 8'd17};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd148, 8'd60, 8'd20};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd136, 8'd53, 8'd3};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd119, 8'd65, 8'd37};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd104, 8'd92, 8'd92};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd99, 8'd121, 8'd135};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd103, 8'd135, 8'd148};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd123, 8'd146, 8'd154};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd164, 8'd173, 8'd180};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd202, 8'd202, 8'd210};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd188, 8'd203, 8'd208};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd157, 8'd193, 8'd189};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd168, 8'd200, 8'd185};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd161, 8'd137, 8'd111};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd178, 8'd79, 8'd38};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd203, 8'd69, 8'd8};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd200, 8'd91, 8'd8};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd181, 8'd113, 8'd14};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd245, 8'd159, 8'd24};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd237, 8'd153, 8'd21};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd229, 8'd145, 8'd21};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd224, 8'd143, 8'd28};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd219, 8'd144, 8'd43};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd212, 8'd141, 8'd53};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd198, 8'd132, 8'd56};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd187, 8'd124, 8'd53};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd193, 8'd130, 8'd61};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd186, 8'd132, 8'd70};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd181, 8'd143, 8'd94};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd186, 8'd168, 8'd132};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd196, 8'd194, 8'd169};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd198, 8'd209, 8'd193};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd188, 8'd208, 8'd197};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd179, 8'd200, 8'd191};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd151, 8'd172, 8'd167};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd124, 8'd146, 8'd143};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd98, 8'd124, 8'd123};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd91, 8'd120, 8'd124};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd98, 8'd133, 8'd139};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd110, 8'd148, 8'd159};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd96, 8'd138, 8'd152};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd66, 8'd109, 8'd125};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd68, 8'd105, 8'd111};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd123, 8'd164, 8'd168};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd131, 8'd176, 8'd179};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd112, 8'd162, 8'd163};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd117, 8'd165, 8'd167};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd123, 8'd167, 8'd170};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd104, 8'd143, 8'd148};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd111, 8'd146, 8'd152};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd76, 8'd101, 8'd98};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd135, 8'd157, 8'd155};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd203, 8'd221, 8'd221};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd165, 8'd184, 8'd190};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd106, 8'd127, 8'd132};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd85, 8'd113, 8'd117};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd96, 8'd129, 8'd134};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd95, 8'd136, 8'd140};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd109, 8'd157, 8'd161};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd129, 8'd180, 8'd183};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd118, 8'd173, 8'd176};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd120, 8'd168, 8'd170};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd138, 8'd183, 8'd186};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd141, 8'd185, 8'd188};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd67, 8'd108, 8'd110};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd89, 8'd129, 8'd129};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd98, 8'd136, 8'd137};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd84, 8'd123, 8'd122};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd88, 8'd127, 8'd126};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd144, 8'd163, 8'd161};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd159, 8'd171, 8'd169};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd176, 8'd181, 8'd175};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd192, 8'd185, 8'd175};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd196, 8'd178, 8'd166};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd190, 8'd161, 8'd145};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd178, 8'd141, 8'd123};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd169, 8'd128, 8'd108};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd166, 8'd102, 8'd64};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd164, 8'd96, 8'd57};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd163, 8'd86, 8'd44};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd162, 8'd78, 8'd32};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd163, 8'd75, 8'd25};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd165, 8'd79, 8'd22};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd169, 8'd85, 8'd25};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd170, 8'd89, 8'd26};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd178, 8'd99, 8'd7};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd201, 8'd118, 8'd22};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd211, 8'd124, 8'd21};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd228, 8'd137, 8'd32};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd215, 8'd119, 8'd17};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd181, 8'd87, 8'd0};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd184, 8'd88, 8'd2};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd180, 8'd84, 8'd7};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd187, 8'd64, 8'd0};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd165, 8'd78, 8'd24};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd139, 8'd102, 8'd83};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd159, 8'd167, 8'd169};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd168, 8'd197, 8'd205};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd163, 8'd194, 8'd199};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd118, 8'd143, 8'd148};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd99, 8'd118, 8'd125};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd108, 8'd103, 8'd97};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd119, 8'd107, 8'd95};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd121, 8'd89, 8'd68};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd122, 8'd59, 8'd28};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd140, 8'd51, 8'd9};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd169, 8'd74, 8'd16};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd189, 8'd110, 8'd35};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd198, 8'd134, 8'd46};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd223, 8'd173, 8'd60};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd226, 8'd187, 8'd70};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd232, 8'd208, 8'd84};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd238, 8'd228, 8'd96};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd247, 8'd241, 8'd105};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd104};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd95};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd253, 8'd221, 8'd86};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd249, 8'd196, 8'd68};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd243, 8'd193, 8'd62};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd48};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd243, 8'd190, 8'd52};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd65};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd247, 8'd180, 8'd49};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd224, 8'd149, 8'd22};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd226, 8'd143, 8'd23};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd245, 8'd164, 8'd49};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd48};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd220, 8'd144, 8'd50};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd217, 8'd147, 8'd61};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd226, 8'd162, 8'd74};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd232, 8'd178, 8'd78};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd234, 8'd187, 8'd73};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd231, 8'd190, 8'd66};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd108};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd101};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd94};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd87};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd88};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd94};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd253, 8'd217, 8'd103};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd108};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd244, 8'd211, 8'd95};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd251, 8'd219, 8'd108};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd254, 8'd227, 8'd124};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd246, 8'd223, 8'd129};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd234, 8'd218, 8'd130};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd233, 8'd221, 8'd135};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd244, 8'd237, 8'd149};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd164};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd251, 8'd224, 8'd153};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd235, 8'd194, 8'd112};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd224, 8'd165, 8'd65};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd234, 8'd157, 8'd39};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd29};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd26};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd252, 8'd175, 8'd19};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd246, 8'd173, 8'd16};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd242, 8'd176, 8'd20};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd245, 8'd168, 8'd12};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd250, 8'd177, 8'd38};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd112};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd253, 8'd245, 8'd199};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd53: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd187};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd239, 8'd202, 8'd114};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd235, 8'd184, 8'd41};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd246, 8'd181, 8'd15};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd23};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd254, 8'd168, 8'd29};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd250, 8'd167, 8'd25};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd24};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd31};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd244, 8'd150, 8'd34};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd233, 8'd156, 8'd52};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd238, 8'd181, 8'd92};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd253, 8'd212, 8'd132};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd156};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd164};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd253, 8'd240, 8'd162};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd254, 8'd229, 8'd126};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd251, 8'd227, 8'd121};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd250, 8'd223, 8'd118};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd248, 8'd220, 8'd113};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd109};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd251, 8'd217, 8'd110};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd254, 8'd217, 8'd111};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd113};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd242, 8'd216, 8'd77};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd244, 8'd215, 8'd87};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd247, 8'd211, 8'd101};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd249, 8'd203, 8'd109};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd249, 8'd195, 8'd109};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd247, 8'd186, 8'd97};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd247, 8'd181, 8'd84};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd75};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd220, 8'd148, 8'd50};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd220, 8'd141, 8'd48};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd229, 8'd141, 8'd52};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd243, 8'd149, 8'd61};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd228, 8'd134, 8'd38};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd214, 8'd126, 8'd16};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd240, 8'd161, 8'd34};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd54};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd75};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd68};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd241, 8'd184, 8'd55};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd228, 8'd179, 8'd51};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd237, 8'd196, 8'd70};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd97};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd108};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd254, 8'd226, 8'd103};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd104};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd248, 8'd219, 8'd101};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd231, 8'd194, 8'd88};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd213, 8'd168, 8'd67};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd195, 8'd141, 8'd43};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd178, 8'd114, 8'd26};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd159, 8'd88, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd148, 8'd70, 8'd22};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd143, 8'd60, 8'd6};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd121, 8'd58, 8'd25};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd109, 8'd78, 8'd73};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd111, 8'd114, 8'd121};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd105, 8'd129, 8'd133};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd102, 8'd128, 8'd127};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd136, 8'd150, 8'd153};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd182, 8'd185, 8'd192};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd199, 8'd217, 8'd219};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd169, 8'd196, 8'd187};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd159, 8'd178, 8'd150};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd141, 8'd113, 8'd65};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd169, 8'd82, 8'd15};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd189, 8'd69, 8'd0};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd196, 8'd90, 8'd6};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd180, 8'd98, 8'd12};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd224, 8'd143, 8'd36};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd223, 8'd141, 8'd33};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd219, 8'd132, 8'd27};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd209, 8'd120, 8'd20};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd196, 8'd108, 8'd19};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd185, 8'd103, 8'd27};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd180, 8'd106, 8'd43};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd179, 8'd110, 8'd53};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd175, 8'd116, 8'd50};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd149, 8'd103, 8'd44};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd117, 8'd90, 8'd45};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd96, 8'd91, 8'd62};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd90, 8'd103, 8'd86};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd91, 8'd116, 8'd110};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd91, 8'd123, 8'd120};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd88, 8'd122, 8'd121};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd102, 8'd133, 8'd128};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd111, 8'd143, 8'd140};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd120, 8'd154, 8'd153};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd120, 8'd155, 8'd157};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd121, 8'd158, 8'd164};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd111, 8'd149, 8'd158};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd92, 8'd132, 8'd142};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd69, 8'd111, 8'd123};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd85, 8'd120, 8'd122};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd117, 8'd157, 8'd157};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd126, 8'd172, 8'd170};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd119, 8'd169, 8'd166};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd119, 8'd169, 8'd166};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd110, 8'd152, 8'd151};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd74, 8'd108, 8'd110};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd82, 8'd111, 8'd115};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd189, 8'd203, 8'd203};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd221, 8'd233, 8'd233};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd227, 8'd238, 8'd240};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd157, 8'd175, 8'd177};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd99, 8'd124, 8'd128};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd95, 8'd129, 8'd131};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd100, 8'd141, 8'd143};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd104, 8'd152, 8'd154};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd127, 8'd176, 8'd180};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd135, 8'd174, 8'd179};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd141, 8'd179, 8'd182};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd117, 8'd150, 8'd155};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd49, 8'd80, 8'd83};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd84, 8'd115, 8'd118};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd109, 8'd143, 8'd144};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd120, 8'd159, 8'd156};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd120, 8'd161, 8'd157};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd94, 8'd128, 8'd129};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd98, 8'd128, 8'd128};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd105, 8'd127, 8'd125};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd112, 8'd124, 8'd120};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd117, 8'd120, 8'd111};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd119, 8'd113, 8'd101};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd120, 8'd106, 8'd93};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd120, 8'd103, 8'd87};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd130, 8'd81, 8'd41};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd136, 8'd78, 8'd38};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd144, 8'd75, 8'd33};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd154, 8'd71, 8'd27};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd158, 8'd67, 8'd22};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd160, 8'd65, 8'd21};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd156, 8'd63, 8'd19};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd154, 8'd63, 8'd18};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd167, 8'd85, 8'd11};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd189, 8'd106, 8'd28};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd202, 8'd116, 8'd31};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd206, 8'd118, 8'd28};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd193, 8'd106, 8'd13};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd177, 8'd92, 8'd0};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd175, 8'd94, 8'd2};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd170, 8'd91, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd184, 8'd73, 8'd0};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd165, 8'd82, 8'd28};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd129, 8'd91, 8'd72};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd131, 8'd135, 8'd136};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd142, 8'd171, 8'd175};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd126, 8'd154, 8'd157};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd95, 8'd106, 8'd110};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd103, 8'd98, 8'd105};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd114, 8'd77, 8'd61};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd122, 8'd84, 8'd61};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd119, 8'd73, 8'd39};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd122, 8'd55, 8'd12};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd143, 8'd57, 8'd6};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd166, 8'd78, 8'd15};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd184, 8'd112, 8'd38};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd200, 8'd144, 8'd61};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd210, 8'd171, 8'd66};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd229, 8'd195, 8'd85};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd246, 8'd221, 8'd103};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd252, 8'd232, 8'd109};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd104};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd96};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd254, 8'd217, 8'd84};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd250, 8'd206, 8'd73};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd239, 8'd183, 8'd48};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd236, 8'd180, 8'd43};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd242, 8'd186, 8'd49};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd66};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd65};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd234, 8'd160, 8'd37};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd214, 8'd130, 8'd16};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd218, 8'd130, 8'd22};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd202, 8'd121, 8'd0};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd217, 8'd137, 8'd14};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd231, 8'd153, 8'd42};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd232, 8'd159, 8'd57};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd226, 8'd157, 8'd62};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd229, 8'd165, 8'd68};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd245, 8'd186, 8'd86};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd99};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd114};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd109};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd100};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd94};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd94};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd98};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd103};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd247, 8'd216, 8'd108};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd253, 8'd230, 8'd124};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd250, 8'd228, 8'd127};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd246, 8'd227, 8'd135};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd247, 8'd229, 8'd143};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd252, 8'd231, 8'd150};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd253, 8'd231, 8'd146};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd251, 8'd226, 8'd136};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd247, 8'd221, 8'd128};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd96};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd226, 8'd168, 8'd71};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd232, 8'd160, 8'd50};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd250, 8'd166, 8'd41};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd29};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd252, 8'd168, 8'd17};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd250, 8'd173, 8'd15};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd25};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd238, 8'd177, 8'd27};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd237, 8'd179, 8'd46};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd245, 8'd200, 8'd99};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd176};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd54: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd249, 8'd228, 8'd181};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd231, 8'd196, 8'd96};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd234, 8'd181, 8'd39};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd247, 8'd182, 8'd20};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd22};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd253, 8'd177, 8'd29};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd250, 8'd175, 8'd34};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd44};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd47};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd246, 8'd156, 8'd44};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd229, 8'd147, 8'd45};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd235, 8'd166, 8'd71};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd114};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd139};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd139};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd147};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd146};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd141};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd134};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd252, 8'd227, 8'd124};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd249, 8'd223, 8'd113};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd245, 8'd220, 8'd102};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd242, 8'd217, 8'd98};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd247, 8'd221, 8'd84};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd248, 8'd217, 8'd92};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd102};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd254, 8'd205, 8'd112};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd253, 8'd199, 8'd113};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd246, 8'd186, 8'd98};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd232, 8'd171, 8'd78};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd222, 8'd160, 8'd61};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd227, 8'd164, 8'd58};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd223, 8'd154, 8'd53};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd227, 8'd146, 8'd54};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd223, 8'd133, 8'd45};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd215, 8'd125, 8'd29};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd207, 8'd121, 8'd12};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd209, 8'd131, 8'd7};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd236, 8'd164, 8'd28};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd253, 8'd191, 8'd56};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd64};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd253, 8'd190, 8'd59};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd235, 8'd174, 8'd47};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd227, 8'd169, 8'd43};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd240, 8'd184, 8'd61};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd82};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd95};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd101};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd241, 8'd213, 8'd103};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd232, 8'd198, 8'd100};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd225, 8'd185, 8'd89};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd216, 8'd168, 8'd70};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd194, 8'd139, 8'd48};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd166, 8'd102, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd145, 8'd76, 8'd19};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd138, 8'd61, 8'd7};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd122, 8'd53, 8'd20};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd115, 8'd68, 8'd58};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd115, 8'd100, 8'd95};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd103, 8'd116, 8'd107};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd89, 8'd115, 8'd102};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd110, 8'd131, 8'd126};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd147, 8'd158, 8'd164};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd181, 8'd199, 8'd211};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd176, 8'd188, 8'd186};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd151, 8'd146, 8'd116};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd145, 8'd107, 8'd44};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd167, 8'd91, 8'd5};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd182, 8'd83, 8'd0};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd191, 8'd88, 8'd9};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd186, 8'd87, 8'd22};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd194, 8'd113, 8'd31};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd212, 8'd123, 8'd39};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd221, 8'd125, 8'd38};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd207, 8'd105, 8'd21};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd178, 8'd76, 8'd1};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd156, 8'd62, 8'd0};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd156, 8'd70, 8'd19};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd165, 8'd86, 8'd43};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd118, 8'd102, 8'd69};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd119, 8'd112, 8'd86};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd119, 8'd127, 8'd112};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd120, 8'd142, 8'd139};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd120, 8'd154, 8'd156};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd123, 8'd161, 8'd164};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd127, 8'd165, 8'd168};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd132, 8'd168, 8'd168};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd123, 8'd164, 8'd160};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd125, 8'd164, 8'd161};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd121, 8'd160, 8'd159};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd116, 8'd154, 8'd155};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd122, 8'd160, 8'd161};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd125, 8'd163, 8'd166};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd119, 8'd154, 8'd160};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd105, 8'd140, 8'd146};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd83, 8'd117, 8'd116};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd109, 8'd148, 8'd145};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd145, 8'd192, 8'd186};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd124, 8'd175, 8'd168};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd102, 8'd151, 8'd145};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd77, 8'd118, 8'd114};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd113, 8'd143, 8'd143};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd195, 8'd216, 8'd219};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd197, 8'd213, 8'd213};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd114, 8'd138, 8'd140};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd84, 8'd115, 8'd117};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd104, 8'd142, 8'd145};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd122, 8'd162, 8'd164};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd138, 8'd178, 8'd178};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd141, 8'd176, 8'd178};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd98, 8'd129, 8'd132};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd77, 8'd107, 8'd109};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd92, 8'd124, 8'd123};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd108, 8'd144, 8'd142};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd112, 8'd155, 8'd148};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd109, 8'd156, 8'd148};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd100, 8'd149, 8'd154};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd105, 8'd153, 8'd157};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd114, 8'd155, 8'd157};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd117, 8'd153, 8'd153};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd113, 8'd142, 8'd138};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd103, 8'd126, 8'd120};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd91, 8'd108, 8'd100};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd82, 8'd98, 8'd88};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd89, 8'd93, 8'd68};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd95, 8'd85, 8'd58};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd106, 8'd73, 8'd40};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd118, 8'd60, 8'd23};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd130, 8'd51, 8'd12};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd139, 8'd46, 8'd5};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd147, 8'd45, 8'd5};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd149, 8'd46, 8'd5};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd167, 8'd76, 8'd5};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd184, 8'd93, 8'd22};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd199, 8'd105, 8'd33};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd184, 8'd90, 8'd16};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd174, 8'd82, 8'd7};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd177, 8'd90, 8'd13};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd166, 8'd85, 8'd6};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd157, 8'd80, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd168, 8'd90, 8'd26};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd138, 8'd78, 8'd41};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd113, 8'd86, 8'd77};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd102, 8'd110, 8'd113};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd106, 8'd131, 8'd128};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd92, 8'd104, 8'd92};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd97, 8'd78, 8'd64};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd118, 8'd69, 8'd62};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd128, 8'd57, 8'd35};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd128, 8'd67, 8'd36};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd122, 8'd63, 8'd19};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd126, 8'd61, 8'd7};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd148, 8'd72, 8'd12};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd164, 8'd85, 8'd19};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd182, 8'd114, 8'd43};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd209, 8'd153, 8'd78};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd223, 8'd188, 8'd96};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd242, 8'd206, 8'd110};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd119};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd112};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd98};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd83};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd242, 8'd184, 8'd58};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd221, 8'd162, 8'd34};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd244, 8'd186, 8'd43};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd244, 8'd186, 8'd43};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd54};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd61};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd238, 8'd169, 8'd42};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd214, 8'd134, 8'd19};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd210, 8'd121, 8'd17};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd216, 8'd122, 8'd26};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd216, 8'd137, 8'd42};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd212, 8'd136, 8'd38};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd211, 8'd138, 8'd36};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd216, 8'd147, 8'd43};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd227, 8'd163, 8'd55};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd241, 8'd181, 8'd67};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd252, 8'd195, 8'd79};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd84};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd210, 8'd89};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd251, 8'd212, 8'd91};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd252, 8'd215, 8'd98};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd254, 8'd218, 8'd104};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd252, 8'd220, 8'd109};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd251, 8'd220, 8'd112};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd248, 8'd219, 8'd115};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd247, 8'd220, 8'd117};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd144};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd249, 8'd229, 8'd143};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd248, 8'd225, 8'd147};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd154};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd154};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd135};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd249, 8'd190, 8'd100};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd233, 8'd167, 8'd71};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd230, 8'd153, 8'd45};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd56};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd58};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd41};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd249, 8'd163, 8'd24};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd20};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd253, 8'd180, 8'd25};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd28};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd240, 8'd181, 8'd43};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd241, 8'd203, 8'd96};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd246, 8'd230, 8'd170};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd254, 8'd252, 8'd229};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd55: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd169};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd236, 8'd192, 8'd71};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd232, 8'd176, 8'd5};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd246, 8'd184, 8'd1};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd253, 8'd184, 8'd29};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd245, 8'd171, 8'd50};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd63};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd59};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd58};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd57};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd249, 8'd158, 8'd51};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd232, 8'd154, 8'd54};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd233, 8'd170, 8'd77};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd243, 8'd192, 8'd103};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd251, 8'd221, 8'd159};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd160};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd158};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd150};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd135};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd251, 8'd232, 8'd114};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd242, 8'd225, 8'd95};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd236, 8'd220, 8'd81};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd254, 8'd211, 8'd116};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd108};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd94};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd81};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd68};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd243, 8'd200, 8'd62};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd230, 8'd185, 8'd58};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd220, 8'd175, 8'd56};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd205, 8'd154, 8'd39};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd209, 8'd148, 8'd41};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd218, 8'd145, 8'd50};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd207, 8'd126, 8'd35};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd214, 8'd130, 8'd34};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd210, 8'd129, 8'd21};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd185, 8'd114, 8'd0};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd201, 8'd135, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd240, 8'd182, 8'd39};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd246, 8'd185, 8'd43};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd54};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd64};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd57};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd242, 8'd173, 8'd46};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd240, 8'd172, 8'd47};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd249, 8'd181, 8'd56};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd249, 8'd227, 8'd108};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd249, 8'd221, 8'd114};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd117};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd239, 8'd198, 8'd106};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd222, 8'd176, 8'd82};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd194, 8'd140, 8'd50};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd160, 8'd101, 8'd25};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd138, 8'd74, 8'd12};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd131, 8'd58, 8'd5};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd123, 8'd53, 8'd19};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd120, 8'd62, 8'd48};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd116, 8'd88, 8'd77};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd99, 8'd103, 8'd86};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd83, 8'd108, 8'd87};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd94, 8'd120, 8'd111};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd118, 8'd136, 8'd140};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd147, 8'd165, 8'd189};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd170, 8'd173, 8'd180};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd145, 8'd124, 8'd97};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd161, 8'd114, 8'd46};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd173, 8'd105, 8'd8};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd187, 8'd100, 8'd5};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd191, 8'd88, 8'd19};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd35};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd172, 8'd85, 8'd16};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd190, 8'd96, 8'd24};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd208, 8'd102, 8'd26};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd204, 8'd92, 8'd16};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd183, 8'd70, 8'd0};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd160, 8'd55, 8'd0};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd149, 8'd54, 8'd10};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd147, 8'd59, 8'd23};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd106, 8'd130, 8'd132};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd117, 8'd148, 8'd153};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd126, 8'd166, 8'd178};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd122, 8'd171, 8'd188};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd112, 8'd161, 8'd178};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd107, 8'd154, 8'd164};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd116, 8'd153, 8'd159};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd127, 8'd159, 8'd158};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd107, 8'd152, 8'd149};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd112, 8'd157, 8'd154};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd112, 8'd154, 8'd152};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd109, 8'd149, 8'd148};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd111, 8'd147, 8'd147};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd123, 8'd157, 8'd158};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd129, 8'd160, 8'd162};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd128, 8'd159, 8'd161};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd114, 8'd144, 8'd142};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd107, 8'd143, 8'd139};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd141, 8'd186, 8'd179};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd104, 8'd155, 8'd146};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd91, 8'd138, 8'd130};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd56, 8'd95, 8'd90};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd135, 8'd161, 8'd160};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd200, 8'd218, 8'd218};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd103, 8'd127, 8'd129};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd76, 8'd106, 8'd108};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd121, 8'd152, 8'd155};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd134, 8'd179, 8'd176};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd138, 8'd178, 8'd177};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd87, 8'd123, 8'd121};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd113, 8'd147, 8'd146};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd109, 8'd145, 8'd141};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd117, 8'd160, 8'd151};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd111, 8'd163, 8'd151};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd114, 8'd170, 8'd157};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd105, 8'd164, 8'd172};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd106, 8'd163, 8'd170};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd109, 8'd164, 8'd169};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd113, 8'd164, 8'd167};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd118, 8'd164, 8'd164};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd123, 8'd165, 8'd163};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd126, 8'd165, 8'd162};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd129, 8'd165, 8'd161};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd122, 8'd175, 8'd165};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd118, 8'd152, 8'd138};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd114, 8'd116, 8'd94};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd114, 8'd79, 8'd49};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd121, 8'd53, 8'd16};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd132, 8'd41, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd145, 8'd40, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd153, 8'd42, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd153, 8'd55, 8'd0};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd169, 8'd71, 8'd0};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd190, 8'd89, 8'd19};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd168, 8'd66, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd164, 8'd66, 8'd3};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd184, 8'd91, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd171, 8'd85, 8'd24};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd162, 8'd81, 8'd18};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd151, 8'd104, 8'd58};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd108, 8'd73, 8'd51};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd97, 8'd85, 8'd87};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd84, 8'd97, 8'd105};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd78, 8'd98, 8'd89};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd72, 8'd68, 8'd43};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd111, 8'd62, 8'd32};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd133, 8'd47, 8'd22};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd142, 8'd52, 8'd26};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd138, 8'd62, 8'd26};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd128, 8'd65, 8'd12};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd133, 8'd72, 8'd9};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd156, 8'd87, 8'd20};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd168, 8'd95, 8'd27};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd185, 8'd120, 8'd52};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd217, 8'd163, 8'd93};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd218, 8'd186, 8'd103};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd248, 8'd210, 8'd125};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd129};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd254, 8'd194, 8'd98};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd235, 8'd166, 8'd62};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd234, 8'd163, 8'd49};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd246, 8'd174, 8'd53};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd253, 8'd184, 8'd57};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd52};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd53};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd61};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd248, 8'd184, 8'd48};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd209, 8'd138, 8'd12};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd197, 8'd115, 8'd5};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd213, 8'd120, 8'd24};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd222, 8'd124, 8'd35};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd201, 8'd131, 8'd43};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd209, 8'd140, 8'd45};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd217, 8'd152, 8'd50};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd221, 8'd161, 8'd51};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd223, 8'd167, 8'd54};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd230, 8'd177, 8'd65};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd244, 8'd192, 8'd83};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd99};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd251, 8'd225, 8'd70};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd222, 8'd76};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd248, 8'd220, 8'd87};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd248, 8'd219, 8'd101};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd249, 8'd221, 8'd114};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd126};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd133};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd137};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd248, 8'd225, 8'd145};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd157};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd164};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd153};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd250, 8'd193, 8'd124};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd241, 8'd168, 8'd91};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd242, 8'd154, 8'd65};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd247, 8'd150, 8'd55};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd48};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd44};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd254, 8'd165, 8'd39};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd251, 8'd167, 8'd35};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd254, 8'd172, 8'd36};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd34};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd252, 8'd181, 8'd27};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd250, 8'd182, 8'd23};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd245, 8'd187, 8'd54};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd249, 8'd222, 8'd133};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd249, 8'd253, 8'd218};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd56: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd227};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd242, 8'd226, 8'd174};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd229, 8'd198, 8'd108};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd233, 8'd180, 8'd52};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd252, 8'd178, 8'd21};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd8};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd250, 8'd180, 8'd58};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd248, 8'd181, 8'd41};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd248, 8'd181, 8'd28};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd253, 8'd184, 8'd31};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd43};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd253, 8'd170, 8'd52};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd243, 8'd155, 8'd45};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd235, 8'd143, 8'd32};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd232, 8'd177, 8'd95};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd244, 8'd191, 8'd113};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd133};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd149};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd150};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd142};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd252, 8'd226, 8'd131};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd250, 8'd226, 8'd126};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd249, 8'd210, 8'd107};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd251, 8'd210, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd253, 8'd211, 8'd99};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd95};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd91};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd250, 8'd197, 8'd81};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd238, 8'd181, 8'd68};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd228, 8'd168, 8'd58};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd226, 8'd158, 8'd57};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd220, 8'd151, 8'd50};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd215, 8'd139, 8'd41};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd213, 8'd130, 8'd34};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd213, 8'd124, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd210, 8'd115, 8'd23};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd204, 8'd105, 8'd14};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd200, 8'd96, 8'd7};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd204, 8'd135, 8'd8};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd248, 8'd181, 8'd48};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd66};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd50};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd249, 8'd189, 8'd43};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd56};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd64};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd64};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd243, 8'd149, 8'd51};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd248, 8'd164, 8'd65};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd253, 8'd183, 8'd85};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd191, 8'd97};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd236, 8'd177, 8'd97};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd209, 8'd144, 8'd80};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd181, 8'd104, 8'd58};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd163, 8'd78, 8'd41};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd135, 8'd63, 8'd15};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd134, 8'd59, 8'd17};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd132, 8'd58, 8'd21};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd126, 8'd59, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd118, 8'd66, 8'd42};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd108, 8'd77, 8'd56};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd97, 8'd89, 8'd66};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd92, 8'd96, 8'd73};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd112, 8'd131, 8'd145};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd130, 8'd146, 8'd143};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd77};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd148, 8'd117, 8'd70};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd182, 8'd117, 8'd61};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd162, 8'd78, 8'd18};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd174, 8'd88, 8'd27};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd161, 8'd81, 8'd20};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd187, 8'd68, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd183, 8'd76, 8'd4};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd186, 8'd93, 8'd26};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd191, 8'd97, 8'd27};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd175, 8'd76, 8'd8};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd140, 8'd57, 8'd5};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd113, 8'd65, 8'd45};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd106, 8'd86, 8'd95};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd127, 8'd149, 8'd147};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd117, 8'd151, 8'd150};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd104, 8'd153, 8'd157};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd96, 8'd157, 8'd162};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd96, 8'd156, 8'd164};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd107, 8'd156, 8'd163};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd122, 8'd152, 8'd160};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd133, 8'd150, 8'd158};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd105, 8'd161, 8'd124};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd96, 8'd132, 8'd118};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd107, 8'd124, 8'd134};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd99, 8'd112, 8'd128};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd107, 8'd132, 8'd137};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd91, 8'd130, 8'd127};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd99, 8'd141, 8'd140};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd115, 8'd155, 8'd163};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd99, 8'd140, 8'd146};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd124, 8'd165, 8'd169};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd131, 8'd173, 8'd172};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd101, 8'd143, 8'd141};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd42, 8'd84, 8'd83};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd77, 8'd118, 8'd122};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd114, 8'd154, 8'd162};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd217, 8'd255, 8'd255};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd230, 8'd243, 8'd249};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd118, 8'd141, 8'd149};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd68, 8'd101, 8'd110};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd93, 8'd133, 8'd143};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd126, 8'd167, 8'd173};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd124, 8'd165, 8'd167};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd104, 8'd145, 8'd141};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd112, 8'd152, 8'd144};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd110, 8'd145, 8'd139};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd110, 8'd138, 8'd139};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd125, 8'd148, 8'd156};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd117, 8'd134, 8'd150};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd116, 8'd141, 8'd135};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd106, 8'd148, 8'd134};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd94, 8'd155, 8'd137};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd94, 8'd158, 8'd141};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd101, 8'd158, 8'd149};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd110, 8'd158, 8'd160};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd111, 8'd161, 8'd170};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd110, 8'd163, 8'd177};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd111, 8'd162, 8'd153};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd125, 8'd175, 8'd176};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd127, 8'd160, 8'd165};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd116, 8'd107, 8'd98};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd116, 8'd57, 8'd25};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd132, 8'd39, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd144, 8'd47, 8'd5};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd143, 8'd54, 8'd24};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd156, 8'd62, 8'd11};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd157, 8'd65, 8'd18};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd144, 8'd55, 8'd11};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd156, 8'd71, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd157, 8'd76, 8'd29};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd144, 8'd67, 8'd11};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd159, 8'd85, 8'd20};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd160, 8'd88, 8'd14};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd134, 8'd97, 8'd71};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd101, 8'd86, 8'd63};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd93, 8'd102, 8'd83};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd90, 8'd104, 8'd89};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd78, 8'd72, 8'd60};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd93, 8'd58, 8'd39};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd119, 8'd64, 8'd33};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd128, 8'd65, 8'd22};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd132, 8'd67, 8'd11};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd138, 8'd71, 8'd18};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd147, 8'd77, 8'd28};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd157, 8'd85, 8'd37};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd170, 8'd97, 8'd46};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd191, 8'd116, 8'd58};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd213, 8'd138, 8'd71};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd230, 8'd153, 8'd81};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd98};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd254, 8'd181, 8'd79};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd58};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd235, 8'd165, 8'd41};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd240, 8'd172, 8'd35};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd248, 8'd183, 8'd39};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd254, 8'd190, 8'd41};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd43};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd254, 8'd197, 8'd46};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd64};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd53};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd215, 8'd125, 8'd15};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd198, 8'd104, 8'd6};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd205, 8'd111, 8'd21};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd202, 8'd114, 8'd25};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd203, 8'd119, 8'd31};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd211, 8'd122, 8'd32};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd215, 8'd127, 8'd37};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd221, 8'd138, 8'd44};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd228, 8'd152, 8'd56};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd236, 8'd167, 8'd66};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd242, 8'd181, 8'd75};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd246, 8'd190, 8'd81};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd248, 8'd194, 8'd85};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd99};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd99};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd101};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd106};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd115};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd247, 8'd218, 8'd126};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd224, 8'd137};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd253, 8'd228, 8'd144};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd142};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd136};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd252, 8'd189, 8'd122};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd241, 8'd166, 8'd99};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd237, 8'd152, 8'd72};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd240, 8'd151, 8'd49};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd251, 8'd162, 8'd34};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd29};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd32};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd250, 8'd168, 8'd32};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd32};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd251, 8'd172, 8'd27};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd249, 8'd183, 8'd24};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd244, 8'd191, 8'd25};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd234, 8'd191, 8'd35};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd225, 8'd187, 8'd44};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd57: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd249, 8'd221, 8'd181};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd243, 8'd202, 8'd112};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd240, 8'd184, 8'd45};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd239, 8'd175, 8'd5};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd249, 8'd182, 8'd7};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd11};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd21};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd37};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd49};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd243, 8'd160, 8'd54};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd52};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd244, 8'd173, 8'd45};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd243, 8'd169, 8'd48};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd237, 8'd166, 8'd52};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd233, 8'd168, 8'd66};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd238, 8'd181, 8'd91};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd250, 8'd202, 8'd120};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd143};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd153};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd154};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd113};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd253, 8'd215, 8'd104};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd249, 8'd210, 8'd93};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd86};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd247, 8'd205, 8'd84};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd246, 8'd200, 8'd80};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd240, 8'd190, 8'd75};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd68};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd225, 8'd150, 8'd49};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd221, 8'd143, 8'd43};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd216, 8'd134, 8'd35};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd216, 8'd127, 8'd33};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd122, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd116, 8'd26};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd212, 8'd106, 8'd18};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd208, 8'd99, 8'd14};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd211, 8'd116, 8'd8};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd221, 8'd135, 8'd16};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd238, 8'd164, 8'd33};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd254, 8'd189, 8'd47};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd49};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd247, 8'd179, 8'd42};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd245, 8'd170, 8'd43};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd55};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd47};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd239, 8'd156, 8'd38};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd223, 8'd148, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd218, 8'd147, 8'd41};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd217, 8'd146, 8'd54};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd210, 8'd137, 8'd60};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd195, 8'd115, 8'd54};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd180, 8'd97, 8'd45};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd158, 8'd74, 8'd28};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd156, 8'd69, 8'd26};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd149, 8'd61, 8'd25};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd138, 8'd55, 8'd25};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd124, 8'd52, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd109, 8'd54, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd96, 8'd58, 8'd37};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd89, 8'd62, 8'd41};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd70, 8'd80, 8'd89};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd72, 8'd87, 8'd84};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd93, 8'd101, 8'd80};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd110, 8'd94, 8'd58};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd138, 8'd87, 8'd42};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd165, 8'd88, 8'd36};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd171, 8'd82, 8'd24};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd176, 8'd86, 8'd23};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd183, 8'd91, 8'd24};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd154, 8'd68, 8'd9};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd147, 8'd62, 8'd8};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd164, 8'd71, 8'd14};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd157, 8'd61, 8'd1};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd129, 8'd48, 8'd1};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd123, 8'd81, 8'd59};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd145, 8'd133, 8'd133};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd121, 8'd155, 8'd157};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd117, 8'd155, 8'd156};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd109, 8'd154, 8'd151};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd102, 8'd147, 8'd142};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd97, 8'd137, 8'd129};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd97, 8'd122, 8'd116};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd99, 8'd108, 8'd105};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd99, 8'd99, 8'd97};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd84, 8'd92, 8'd55};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd94, 8'd88, 8'd66};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd95, 8'd76, 8'd70};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd97, 8'd78, 8'd72};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd92, 8'd90, 8'd77};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd92, 8'd109, 8'd91};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd78, 8'd108, 8'd100};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd53, 8'd86, 8'd91};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd70, 8'd111, 8'd117};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd95, 8'd136, 8'd140};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd111, 8'd152, 8'd154};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd97, 8'd139, 8'd138};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd47, 8'd88, 8'd90};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd68, 8'd109, 8'd115};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd87, 8'd127, 8'd137};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd176, 8'd215, 8'd230};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd198, 8'd213, 8'd220};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd100, 8'd127, 8'd138};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd64, 8'd102, 8'd113};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd55, 8'd99, 8'd112};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd112, 8'd147, 8'd149};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd107, 8'd147, 8'd147};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd101, 8'd145, 8'd146};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd118, 8'd162, 8'd161};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd98, 8'd137, 8'd136};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd80, 8'd106, 8'd107};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd82, 8'd93, 8'd97};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd98, 8'd99, 8'd104};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd110, 8'd94, 8'd94};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd103, 8'd102, 8'd97};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd103};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd102, 8'd124, 8'd111};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd111, 8'd132, 8'd125};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd116, 8'd142, 8'd141};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd113, 8'd153, 8'd153};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd109, 8'd160, 8'd161};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd95, 8'd143, 8'd147};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd98, 8'd152, 8'd164};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd104, 8'd152, 8'd166};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd111, 8'd127, 8'd126};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd122, 8'd88, 8'd61};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd132, 8'd55, 8'd11};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd139, 8'd41, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd143, 8'd40, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd146, 8'd53, 8'd10};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd144, 8'd53, 8'd9};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd132, 8'd43, 8'd0};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd141, 8'd54, 8'd9};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd151, 8'd71, 8'd22};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd145, 8'd69, 8'd19};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd145, 8'd76, 8'd21};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd148, 8'd82, 8'd24};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd126, 8'd99, 8'd80};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd121, 8'd113, 8'd94};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd86, 8'd97, 8'd81};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd90, 8'd98, 8'd85};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd108, 8'd92, 8'd77};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd117, 8'd70, 8'd50};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd137, 8'd71, 8'd37};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd131, 8'd57, 8'd12};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd163, 8'd88, 8'd31};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd168, 8'd93, 8'd38};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd175, 8'd98, 8'd44};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd182, 8'd103, 8'd47};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd190, 8'd110, 8'd49};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd202, 8'd122, 8'd53};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd219, 8'd137, 8'd61};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd230, 8'd149, 8'd67};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd221, 8'd142, 8'd39};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd231, 8'd153, 8'd45};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd48};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd248, 8'd175, 8'd46};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd248, 8'd176, 8'd38};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd248, 8'd177, 8'd35};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd250, 8'd182, 8'd39};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd254, 8'd186, 8'd41};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd250, 8'd178, 8'd42};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd245, 8'd166, 8'd39};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd225, 8'd134, 8'd20};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd206, 8'd107, 8'd6};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd215, 8'd112, 8'd20};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd219, 8'd119, 8'd31};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd206, 8'd112, 8'd24};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd200, 8'd111, 8'd21};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd208, 8'd120, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd213, 8'd128, 8'd35};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd221, 8'd141, 8'd46};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd232, 8'd158, 8'd59};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd243, 8'd176, 8'd72};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd252, 8'd191, 8'd84};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd91};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd96};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd96};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd218, 8'd97};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd251, 8'd216, 8'd100};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd251, 8'd213, 8'd104};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd254, 8'd212, 8'd110};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd116};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd121};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd124};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd237, 8'd171, 8'd84};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd235, 8'd167, 8'd70};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd235, 8'd164, 8'd50};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd243, 8'd169, 8'd38};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd253, 8'd176, 8'd36};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd38};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd250, 8'd172, 8'd36};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd34};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd46};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd43};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd249, 8'd187, 8'd6};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd230, 8'd179, 8'd0};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd226, 8'd185, 8'd43};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd244, 8'd206, 8'd121};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd187};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd58: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd185};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd238, 8'd208, 8'd120};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd222, 8'd189, 8'd74};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd235, 8'd174, 8'd0};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd248, 8'd179, 8'd0};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd7};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd24};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd41};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd252, 8'd168, 8'd52};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd246, 8'd175, 8'd57};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd242, 8'd183, 8'd55};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd26};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd251, 8'd160, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd38};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd234, 8'd157, 8'd49};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd231, 8'd165, 8'd68};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd236, 8'd179, 8'd89};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd246, 8'd196, 8'd109};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd253, 8'd209, 8'd122};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd106};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd101};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd94};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd89};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd86};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd247, 8'd203, 8'd78};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd235, 8'd191, 8'd70};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd225, 8'd180, 8'd61};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd236, 8'd157, 8'd56};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd231, 8'd149, 8'd49};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd224, 8'd138, 8'd39};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd219, 8'd129, 8'd33};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd219, 8'd121, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd215, 8'd111, 8'd22};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd209, 8'd100, 8'd15};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd202, 8'd92, 8'd7};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd205, 8'd89, 8'd2};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd202, 8'd95, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd220, 8'd129, 8'd14};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd251, 8'd174, 8'd44};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd50};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd38};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd247, 8'd178, 8'd39};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd55};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd40};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd253, 8'd171, 8'd33};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd242, 8'd158, 8'd26};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd230, 8'd141, 8'd21};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd217, 8'd126, 8'd21};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd199, 8'd111, 8'd21};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd181, 8'd98, 8'd20};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd171, 8'd89, 8'd16};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd171, 8'd77, 8'd26};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd169, 8'd72, 8'd27};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd167, 8'd65, 8'd25};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd162, 8'd59, 8'd28};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd153, 8'd55, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd141, 8'd55, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd133, 8'd57, 8'd34};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd127, 8'd59, 8'd36};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd73, 8'd67, 8'd67};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd68, 8'd77, 8'd72};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd87, 8'd105, 8'd93};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd92, 8'd95, 8'd76};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd110, 8'd80, 8'd54};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd150, 8'd82, 8'd43};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd170, 8'd76, 8'd24};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd181, 8'd77, 8'd14};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd141, 8'd79, 8'd28};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd119, 8'd52, 8'd7};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd120, 8'd43, 8'd1};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd145, 8'd53, 8'd12};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd144, 8'd55, 8'd11};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd120, 8'd54, 8'd19};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd114, 8'd89, 8'd69};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd131, 8'd137, 8'd133};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd108, 8'd148, 8'd158};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd105, 8'd140, 8'd142};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd103, 8'd126, 8'd116};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd98, 8'd110, 8'd88};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd99, 8'd95, 8'd68};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd100, 8'd83, 8'd57};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd104, 8'd76, 8'd54};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd107, 8'd72, 8'd53};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd126, 8'd70, 8'd33};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd151, 8'd87, 8'd59};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd140, 8'd74, 8'd48};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd151, 8'd92, 8'd60};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd141, 8'd102, 8'd63};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd163, 8'd152, 8'd120};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd147, 8'd161, 8'd148};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd80, 8'd109, 8'd113};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd49, 8'd92, 8'd99};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd63, 8'd106, 8'd112};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd80, 8'd124, 8'd127};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd82, 8'd126, 8'd127};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd47, 8'd91, 8'd94};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd53, 8'd96, 8'd103};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd59, 8'd101, 8'd113};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd134, 8'd176, 8'd192};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd155, 8'd175, 8'd186};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd72, 8'd105, 8'd120};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd56, 8'd99, 8'd115};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd28, 8'd79, 8'd96};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd113, 8'd142, 8'd138};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd112, 8'd150, 8'd151};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd77, 8'd126, 8'd131};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd49, 8'd102, 8'd110};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd58, 8'd101, 8'd107};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd124, 8'd142, 8'd142};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd123, 8'd116, 8'd108};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd110, 8'd83, 8'd72};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd121, 8'd60, 8'd57};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd117, 8'd67, 8'd58};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd117, 8'd75, 8'd61};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd119, 8'd83, 8'd67};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd122, 8'd90, 8'd75};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd116, 8'd100, 8'd85};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd101, 8'd112, 8'd95};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd88, 8'd121, 8'd100};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd95, 8'd125, 8'd133};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd91, 8'd139, 8'd153};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd101, 8'd160, 8'd176};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd117, 8'd165, 8'd169};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd127, 8'd131, 8'd114};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd127, 8'd79, 8'd39};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd135, 8'd45, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd148, 8'd37, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd130, 8'd40, 8'd6};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd128, 8'd36, 8'd0};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd129, 8'd38, 8'd0};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd134, 8'd48, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd148, 8'd68, 8'd17};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd137, 8'd66, 8'd22};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd119, 8'd57, 8'd20};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd134, 8'd78, 8'd45};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd154, 8'd144, 8'd135};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd155, 8'd155, 8'd145};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd77};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd75, 8'd69, 8'd57};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd114, 8'd78, 8'd62};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd134, 8'd68, 8'd42};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd163, 8'd78, 8'd39};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd157, 8'd67, 8'd17};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd174, 8'd85, 8'd25};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd181, 8'd92, 8'd32};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd190, 8'd100, 8'd38};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd196, 8'd107, 8'd39};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd201, 8'd111, 8'd35};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd208, 8'd118, 8'd32};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd217, 8'd128, 8'd34};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd225, 8'd137, 8'd37};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd235, 8'd150, 8'd33};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd243, 8'd159, 8'd37};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd251, 8'd169, 8'd41};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd254, 8'd173, 8'd40};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd252, 8'd175, 8'd37};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd252, 8'd176, 8'd38};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd45};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd52};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd56};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd235, 8'd143, 8'd34};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd199, 8'd97, 8'd0};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd190, 8'd82, 8'd0};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd206, 8'd97, 8'd12};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd211, 8'd107, 8'd20};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd206, 8'd111, 8'd21};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd207, 8'd118, 8'd24};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd221, 8'd138, 8'd44};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd220, 8'd140, 8'd43};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd221, 8'd146, 8'd45};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd226, 8'd155, 8'd51};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd232, 8'd168, 8'd60};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd241, 8'd184, 8'd69};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd250, 8'd198, 8'd80};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd87};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd232, 8'd209, 8'd81};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd242, 8'd214, 8'd89};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd98};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd104};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd99};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd86};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd244, 8'd173, 8'd69};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd234, 8'd159, 8'd57};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd237, 8'd150, 8'd44};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd242, 8'd156, 8'd37};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd250, 8'd164, 8'd29};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd23};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd254, 8'd175, 8'd20};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd250, 8'd177, 8'd23};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd246, 8'd178, 8'd33};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd245, 8'd178, 8'd38};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd29};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd251, 8'd188, 8'd25};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd239, 8'd190, 8'd25};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd232, 8'd197, 8'd55};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd238, 8'd212, 8'd125};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd218};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd59: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd231, 8'd189, 8'd87};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd234, 8'd184, 8'd53};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd243, 8'd178, 8'd14};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd0};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd10};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd253, 8'd179, 8'd46};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd242, 8'd177, 8'd49};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd45};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd48};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd46};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd249, 8'd163, 8'd42};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd238, 8'd155, 8'd33};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd234, 8'd154, 8'd29};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd236, 8'd161, 8'd34};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd242, 8'd169, 8'd41};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd254, 8'd191, 8'd77};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd76};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd74};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd76};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd79};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd76};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd246, 8'd190, 8'd69};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd236, 8'd181, 8'd62};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd233, 8'd159, 8'd52};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd228, 8'd151, 8'd45};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd222, 8'd140, 8'd38};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd219, 8'd133, 8'd34};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd217, 8'd127, 8'd31};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd214, 8'd119, 8'd27};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd209, 8'd109, 8'd21};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd203, 8'd102, 8'd14};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd216, 8'd100, 8'd25};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd189, 8'd83, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd181, 8'd88, 8'd0};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd204, 8'd124, 8'd3};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd238, 8'd164, 8'd31};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd52};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd48};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd254, 8'd171, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd249, 8'd178, 8'd28};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd241, 8'd135, 8'd25};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd217, 8'd117, 8'd21};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd194, 8'd102, 8'd15};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd180, 8'd95, 8'd14};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd161, 8'd67, 8'd5};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd162, 8'd63, 8'd6};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd163, 8'd59, 8'd8};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd161, 8'd54, 8'd10};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd159, 8'd51, 8'd13};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd154, 8'd49, 8'd17};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd149, 8'd50, 8'd19};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd145, 8'd50, 8'd20};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd104, 8'd74, 8'd64};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd104, 8'd100, 8'd91};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd73, 8'd94, 8'd89};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd95, 8'd115, 8'd113};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd123, 8'd112, 8'd106};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd125, 8'd71, 8'd47};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd155, 8'd64, 8'd19};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd167, 8'd57, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd138, 8'd82, 8'd33};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd136, 8'd69, 8'd24};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd131, 8'd48, 8'd8};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd124, 8'd31, 8'd0};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd117, 8'd37, 8'd10};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd111, 8'd68, 8'd49};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd104, 8'd107, 8'd98};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd98, 8'd132, 8'd131};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd71, 8'd98, 8'd109};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd77, 8'd89, 8'd87};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd84, 8'd76, 8'd55};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd96, 8'd62, 8'd25};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd110, 8'd56, 8'd10};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd122, 8'd55, 8'd10};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd133, 8'd59, 8'd20};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd138, 8'd63, 8'd31};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd141, 8'd38, 8'd5};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd157, 8'd57, 8'd23};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd140, 8'd42, 8'd3};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd145, 8'd57, 8'd9};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd134, 8'd67, 8'd15};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd158, 8'd124, 8'd86};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd160, 8'd166, 8'd154};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd84, 8'd117, 8'd126};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd54, 8'd97, 8'd106};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd51, 8'd94, 8'd101};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd54, 8'd97, 8'd103};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd61, 8'd105, 8'd108};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd42, 8'd85, 8'd91};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd41, 8'd84, 8'd93};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd47, 8'd89, 8'd103};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd110, 8'd151, 8'd169};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd223, 8'd236, 8'd244};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd113, 8'd141, 8'd155};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd50, 8'd88, 8'd107};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd43, 8'd91, 8'd111};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd35, 8'd90, 8'd110};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd104, 8'd127, 8'd121};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd73, 8'd108, 8'd110};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd36, 8'd88, 8'd99};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd45, 8'd103, 8'd117};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd93, 8'd136, 8'd145};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd165, 8'd174, 8'd171};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd139, 8'd111, 8'd90};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd127, 8'd72, 8'd42};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd142, 8'd61, 8'd34};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd141, 8'd65, 8'd33};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd145, 8'd69, 8'd35};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd152, 8'd72, 8'd35};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd155, 8'd75, 8'd38};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd144, 8'd82, 8'd43};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd123, 8'd92, 8'd46};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd106, 8'd100, 8'd48};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd105, 8'd99, 8'd87};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd85, 8'd104, 8'd100};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd74, 8'd125, 8'd126};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd84, 8'd146, 8'd145};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd100, 8'd138, 8'd125};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd109, 8'd100, 8'd69};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd124, 8'd61, 8'd17};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd139, 8'd42, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd125, 8'd36, 8'd6};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd123, 8'd33, 8'd0};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd141, 8'd50, 8'd3};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd144, 8'd57, 8'd4};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd141, 8'd63, 8'd14};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd115, 8'd49, 8'd14};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd95, 8'd43, 8'd22};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd137, 8'd93, 8'd84};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd167, 8'd168, 8'd170};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd153, 8'd159, 8'd155};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd102, 8'd103, 8'd95};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd98, 8'd75, 8'd61};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd130, 8'd72, 8'd52};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd151, 8'd62, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd165, 8'd63, 8'd15};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd158, 8'd53, 8'd0};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd172, 8'd70, 8'd4};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd182, 8'd81, 8'd11};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd196, 8'd96, 8'd20};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd206, 8'd107, 8'd22};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd214, 8'd115, 8'd21};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd220, 8'd123, 8'd18};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd227, 8'd131, 8'd18};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd233, 8'd138, 8'd20};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd249, 8'd160, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd248, 8'd160, 8'd27};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd250, 8'd164, 8'd27};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd34};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd43};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd47};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd48};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd249, 8'd170, 8'd43};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd194, 8'd108, 8'd5};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd196, 8'd106, 8'd9};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd186, 8'd87, 8'd0};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd196, 8'd92, 8'd7};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd212, 8'd108, 8'd23};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd208, 8'd110, 8'd21};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd206, 8'd117, 8'd23};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd207, 8'd125, 8'd26};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd210, 8'd128, 8'd29};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd213, 8'd133, 8'd34};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd221, 8'd144, 8'd40};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd229, 8'd158, 8'd50};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd240, 8'd174, 8'd61};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd249, 8'd189, 8'd69};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd77};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd81};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd198, 8'd76};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd247, 8'd193, 8'd71};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd244, 8'd184, 8'd62};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd240, 8'd174, 8'd52};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd240, 8'd166, 8'd45};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd240, 8'd159, 8'd41};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd242, 8'd156, 8'd37};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd244, 8'd155, 8'd37};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd251, 8'd167, 8'd35};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd45};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd55};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd56};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd47};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd252, 8'd172, 8'd35};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd252, 8'd181, 8'd27};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd254, 8'd189, 8'd25};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd237, 8'd176, 8'd0};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd234, 8'd174, 8'd15};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd235, 8'd180, 8'd64};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd242, 8'd199, 8'd120};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd175};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd220};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd60: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd246, 8'd235, 8'd207};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd239, 8'd218, 8'd153};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd235, 8'd195, 8'd84};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd237, 8'd176, 8'd33};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd244, 8'd170, 8'd13};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd251, 8'd171, 8'd14};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd253, 8'd175, 8'd17};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd252, 8'd178, 8'd17};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd253, 8'd181, 8'd45};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd249, 8'd176, 8'd38};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd250, 8'd170, 8'd33};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd32};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd32};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd22};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd254, 8'd145, 8'd14};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd245, 8'd158, 8'd42};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd241, 8'd156, 8'd37};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd240, 8'd156, 8'd32};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd245, 8'd163, 8'd37};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd252, 8'd172, 8'd47};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd57};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd64};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd66};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd241, 8'd171, 8'd59};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd234, 8'd162, 8'd51};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd224, 8'd150, 8'd43};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd218, 8'd139, 8'd36};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd214, 8'd130, 8'd32};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd207, 8'd120, 8'd25};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd198, 8'd107, 8'd16};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd190, 8'd99, 8'd10};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd191, 8'd94, 8'd17};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd186, 8'd94, 8'd9};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd191, 8'd107, 8'd8};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd193, 8'd116, 8'd2};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd198, 8'd120, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd226, 8'd144, 8'd9};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd26};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd46};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd36};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd251, 8'd157, 8'd25};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd253, 8'd147, 8'd27};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd254, 8'd144, 8'd33};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd243, 8'd137, 8'd37};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd219, 8'd121, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd200, 8'd108, 8'd21};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd180, 8'd89, 8'd10};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd178, 8'd85, 8'd8};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd175, 8'd76, 8'd8};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd169, 8'd67, 8'd5};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd161, 8'd55, 8'd3};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd152, 8'd45, 8'd0};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd144, 8'd38, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd138, 8'd34, 8'd0};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd113, 8'd54, 8'd36};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd105, 8'd78, 8'd67};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd60, 8'd74, 8'd74};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd96, 8'd123, 8'd130};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd152, 8'd155, 8'd160};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd128, 8'd88, 8'd78};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd118, 8'd38, 8'd5};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd143, 8'd39, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd145, 8'd74, 8'd20};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd167, 8'd81, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd169, 8'd71, 8'd24};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd145, 8'd48, 8'd13};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd120, 8'd54, 8'd32};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd109, 8'd87, 8'd76};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd88, 8'd109, 8'd104};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd61, 8'd110, 8'd107};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd79, 8'd74, 8'd71};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd92, 8'd73, 8'd59};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd115, 8'd70, 8'd39};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd139, 8'd69, 8'd20};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd157, 8'd68, 8'd10};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd168, 8'd69, 8'd10};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd171, 8'd70, 8'd18};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd173, 8'd71, 8'd23};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd167, 8'd55, 8'd18};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd166, 8'd60, 8'd21};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd150, 8'd49, 8'd3};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd144, 8'd47, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd135, 8'd49, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd130, 8'd80, 8'd45};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd151, 8'd151, 8'd143};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd92, 8'd130, 8'd141};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd59, 8'd103, 8'd116};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd46, 8'd90, 8'd101};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd38, 8'd83, 8'd89};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd44, 8'd89, 8'd95};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd37, 8'd82, 8'd88};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd30, 8'd74, 8'd85};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd36, 8'd79, 8'd96};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd85, 8'd128, 8'd147};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd172, 8'd197, 8'd204};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd190, 8'd212, 8'd225};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd72, 8'd107, 8'd126};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd40, 8'd85, 8'd106};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd30, 8'd82, 8'd103};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd44, 8'd101, 8'd120};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd59, 8'd85, 8'd82};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd49, 8'd88, 8'd93};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd41, 8'd95, 8'd107};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd57, 8'd113, 8'd128};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd107, 8'd142, 8'd148};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd158, 8'd151, 8'd141};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd128, 8'd79, 8'd49};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd121, 8'd42, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd143, 8'd66, 8'd10};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd149, 8'd73, 8'd15};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd164, 8'd83, 8'd20};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd184, 8'd90, 8'd26};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd201, 8'd99, 8'd35};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd202, 8'd109, 8'd42};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd189, 8'd121, 8'd46};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd176, 8'd131, 8'd50};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd153, 8'd109, 8'd62};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd116, 8'd97, 8'd57};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd73, 8'd93, 8'd65};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd57, 8'd106, 8'd87};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd71, 8'd119, 8'd105};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd102, 8'd117, 8'd94};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd133, 8'd99, 8'd62};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd153, 8'd83, 8'd34};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd144, 8'd61, 8'd21};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd139, 8'd52, 8'd7};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd157, 8'd65, 8'd16};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd151, 8'd61, 8'd11};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd124, 8'd45, 8'd4};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd91, 8'd31, 8'd5};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd94, 8'd54, 8'd46};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd159, 8'd133, 8'd136};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd165, 8'd176, 8'd180};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd124, 8'd130, 8'd128};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd118, 8'd108, 8'd98};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd118, 8'd75, 8'd56};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd131, 8'd50, 8'd21};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd163, 8'd56, 8'd14};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd172, 8'd59, 8'd1};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd178, 8'd69, 8'd0};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd191, 8'd81, 8'd4};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd203, 8'd94, 8'd12};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd216, 8'd111, 8'd19};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd228, 8'd125, 8'd24};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd236, 8'd134, 8'd23};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd242, 8'd142, 8'd22};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd248, 8'd149, 8'd22};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd253, 8'd156, 8'd25};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd247, 8'd157, 8'd17};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd249, 8'd162, 8'd21};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd254, 8'd169, 8'd27};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd34};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd37};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd239, 8'd162, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd214, 8'd139, 8'd12};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd197, 8'd121, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd186, 8'd110, 8'd12};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd200, 8'd120, 8'd25};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd187, 8'd97, 8'd9};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd190, 8'd94, 8'd10};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd200, 8'd104, 8'd18};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd198, 8'd107, 8'd16};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd205, 8'd123, 8'd24};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd203, 8'd125, 8'd24};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd219, 8'd131, 8'd33};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd226, 8'd140, 8'd39};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd236, 8'd153, 8'd47};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd244, 8'd166, 8'd55};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd250, 8'd175, 8'd58};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd250, 8'd180, 8'd58};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd247, 8'd179, 8'd52};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd243, 8'd178, 8'd48};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd252, 8'd155, 8'd42};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd247, 8'd150, 8'd37};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd240, 8'd145, 8'd27};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd236, 8'd144, 8'd21};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd239, 8'd147, 8'd22};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd245, 8'd156, 8'd26};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd34};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd40};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd250, 8'd179, 8'd35};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd247, 8'd174, 8'd35};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd249, 8'd171, 8'd37};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd44};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd45};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd39};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd25};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd245, 8'd178, 8'd12};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd221, 8'd178, 8'd11};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd234, 8'd192, 8'd71};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd253, 8'd213, 8'd154};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd220};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd61: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd253, 8'd251, 8'd228};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd251, 8'd232, 8'd189};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd243, 8'd205, 8'd142};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd235, 8'd181, 8'd95};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd235, 8'd170, 8'd54};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd173, 8'd17};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd249, 8'd181, 8'd0};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd246, 8'd193, 8'd25};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd247, 8'd190, 8'd25};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd249, 8'd183, 8'd24};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd26};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd31};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd37};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd43};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd45};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd246, 8'd150, 8'd29};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd242, 8'd146, 8'd23};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd239, 8'd144, 8'd18};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd241, 8'd146, 8'd18};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd247, 8'd149, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd249, 8'd150, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd247, 8'd148, 8'd31};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd244, 8'd144, 8'd32};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd234, 8'd157, 8'd43};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd227, 8'd149, 8'd38};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd221, 8'd140, 8'd32};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd217, 8'd131, 8'd28};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd214, 8'd126, 8'd28};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd209, 8'd118, 8'd25};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd202, 8'd108, 8'd20};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd196, 8'd100, 8'd14};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd174, 8'd82, 8'd0};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd189, 8'd104, 8'd13};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd232, 8'd154, 8'd54};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd247, 8'd175, 8'd65};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd212, 8'd142, 8'd21};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd201, 8'd123, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd229, 8'd144, 8'd15};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd254, 8'd163, 8'd31};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd48};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd251, 8'd175, 8'd40};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd246, 8'd162, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd247, 8'd153, 8'd27};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd248, 8'd149, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd243, 8'd143, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd232, 8'd133, 8'd29};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd224, 8'd124, 8'd26};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd212, 8'd116, 8'd16};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd208, 8'd111, 8'd16};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd200, 8'd102, 8'd15};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd189, 8'd89, 8'd11};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd176, 8'd75, 8'd7};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd162, 8'd59, 8'd1};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd150, 8'd46, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd142, 8'd40, 8'd0};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd131, 8'd41, 8'd17};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd98, 8'd46, 8'd32};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd88, 8'd84, 8'd81};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd104, 8'd124, 8'd131};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd167, 8'd176, 8'd185};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd164, 8'd136, 8'd133};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd93, 8'd31, 8'd10};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd114, 8'd30, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd128, 8'd45, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd158, 8'd59, 8'd4};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd180, 8'd71, 8'd15};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd171, 8'd74, 8'd29};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd139, 8'd78, 8'd49};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd106, 8'd85, 8'd66};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd77, 8'd88, 8'd71};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd63, 8'd86, 8'd66};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd141, 8'd105, 8'd73};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd149, 8'd104, 8'd65};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd164, 8'd102, 8'd53};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd178, 8'd99, 8'd40};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd189, 8'd97, 8'd32};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd193, 8'd96, 8'd28};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd192, 8'd94, 8'd29};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd192, 8'd94, 8'd31};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd174, 8'd80, 8'd29};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd160, 8'd74, 8'd23};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd156, 8'd70, 8'd19};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd154, 8'd58, 8'd8};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd150, 8'd53, 8'd8};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd126, 8'd59, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd144, 8'd134, 8'd124};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd114, 8'd152, 8'd155};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd60, 8'd103, 8'd119};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd50, 8'd94, 8'd107};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd40, 8'd84, 8'd95};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd43, 8'd87, 8'd96};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd43, 8'd87, 8'd98};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd28, 8'd71, 8'd87};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd29, 8'd72, 8'd91};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd58, 8'd100, 8'd122};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd114, 8'd148, 8'd157};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd194, 8'd221, 8'd228};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd219, 8'd238, 8'd245};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd143, 8'd172, 8'd188};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd44, 8'd82, 8'd103};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd42, 8'd89, 8'd109};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd29, 8'd80, 8'd99};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd41, 8'd94, 8'd110};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd37, 8'd74, 8'd80};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd56, 8'd100, 8'd109};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd58, 8'd110, 8'd123};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd54, 8'd101, 8'd111};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd105, 8'd125, 8'd124};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd145, 8'd122, 8'd104};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd141, 8'd76, 8'd38};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd137, 8'd42, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd138, 8'd67, 8'd1};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd147, 8'd79, 8'd8};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd164, 8'd95, 8'd17};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd192, 8'd111, 8'd29};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd218, 8'd126, 8'd41};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd230, 8'd140, 8'd52};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd228, 8'd153, 8'd60};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd220, 8'd162, 8'd63};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd222, 8'd160, 8'd83};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd196, 8'd150, 8'd75};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd149, 8'd133, 8'd71};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd100, 8'd115, 8'd72};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd72, 8'd102, 8'd74};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd87, 8'd102, 8'd73};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd136, 8'd114, 8'd73};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd182, 8'd129, 8'd75};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd174, 8'd98, 8'd40};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd164, 8'd79, 8'd24};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd161, 8'd69, 8'd20};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd141, 8'd48, 8'd7};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd102, 8'd22, 8'd0};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd88, 8'd35, 8'd19};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd123, 8'd95, 8'd92};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd180, 8'd169, 8'd173};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd149, 8'd158, 8'd163};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd98, 8'd99, 8'd94};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd120, 8'd94, 8'd79};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd125, 8'd61, 8'd34};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd132, 8'd33, 8'd0};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd177, 8'd57, 8'd4};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd189, 8'd75, 8'd5};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd211, 8'd106, 8'd25};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd216, 8'd107, 8'd16};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd225, 8'd117, 8'd19};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd237, 8'd131, 8'd22};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd244, 8'd141, 8'd23};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd246, 8'd147, 8'd18};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd249, 8'd151, 8'd18};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd253, 8'd157, 8'd21};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd23};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd28};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd29};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd29};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd241, 8'd166, 8'd23};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd227, 8'd156, 8'd16};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd216, 8'd148, 8'd15};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd215, 8'd147, 8'd22};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd215, 8'd149, 8'd27};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd254, 8'd185, 8'd84};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd247, 8'd171, 8'd77};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd199, 8'd111, 8'd22};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd188, 8'd92, 8'd8};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd200, 8'd100, 8'd15};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd201, 8'd106, 8'd16};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd217, 8'd127, 8'd31};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd211, 8'd128, 8'd26};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd241, 8'd143, 8'd44};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd239, 8'd141, 8'd40};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd235, 8'd140, 8'd34};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd230, 8'd138, 8'd27};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd226, 8'd140, 8'd21};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd226, 8'd142, 8'd17};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd226, 8'd145, 8'd14};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd227, 8'd146, 8'd13};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd249, 8'd132, 8'd19};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd253, 8'd138, 8'd23};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd148, 8'd29};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd32};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd34};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd31};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd28};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd248, 8'd172, 8'd26};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd249, 8'd184, 8'd38};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd245, 8'd180, 8'd24};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd241, 8'd178, 8'd5};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd0};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd238, 8'd178, 8'd2};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd239, 8'd180, 8'd24};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd239, 8'd182, 8'd49};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd238, 8'd183, 8'd66};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd240, 8'd214, 8'd130};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd174};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd226};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd62: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd248, 8'd223, 8'd192};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd242, 8'd204, 8'd142};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd241, 8'd193, 8'd91};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd243, 8'd191, 8'd56};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd245, 8'd186, 8'd34};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd251, 8'd190, 8'd37};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd37};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd254, 8'd185, 8'd32};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd249, 8'd173, 8'd27};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd248, 8'd166, 8'd28};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd39};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd50};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd37};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd254, 8'd163, 8'd31};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd160, 8'd27};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd253, 8'd156, 8'd23};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd252, 8'd153, 8'd23};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd247, 8'd145, 8'd21};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd237, 8'd132, 8'd14};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd228, 8'd123, 8'd8};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd216, 8'd118, 8'd9};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd213, 8'd115, 8'd8};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd212, 8'd111, 8'd7};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd216, 8'd112, 8'd15};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd223, 8'd115, 8'd24};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd227, 8'd117, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd225, 8'd113, 8'd31};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd222, 8'd109, 8'd29};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd209, 8'd103, 8'd15};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd191, 8'd94, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd222, 8'd140, 8'd40};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd88};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd82};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd240, 8'd185, 8'd59};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd237, 8'd180, 8'd51};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd228, 8'd169, 8'd39};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd239, 8'd165, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd31};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd244, 8'd173, 8'd31};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd244, 8'd172, 8'd28};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd244, 8'd164, 8'd25};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd244, 8'd156, 8'd22};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd248, 8'd150, 8'd25};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd252, 8'd148, 8'd27};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd231, 8'd117, 8'd5};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd226, 8'd113, 8'd7};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd216, 8'd106, 8'd8};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd205, 8'd97, 8'd9};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd189, 8'd83, 8'd9};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd172, 8'd68, 8'd5};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd160, 8'd55, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd153, 8'd47, 8'd0};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd156, 8'd37, 8'd13};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd121, 8'd46, 8'd27};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd118, 8'd95, 8'd87};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd105, 8'd115, 8'd117};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd149, 8'd156, 8'd164};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd186, 8'd167, 8'd169};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd125, 8'd78, 8'd68};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd95, 8'd35, 8'd11};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd122, 8'd37, 8'd6};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd140, 8'd42, 8'd0};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd161, 8'd55, 8'd0};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd162, 8'd69, 8'd12};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd137, 8'd75, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd115, 8'd80, 8'd40};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd123, 8'd96, 8'd49};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd145, 8'd116, 8'd60};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd192, 8'd135, 8'd68};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd192, 8'd135, 8'd68};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd193, 8'd132, 8'd65};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd194, 8'd131, 8'd62};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd194, 8'd130, 8'd58};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd195, 8'd127, 8'd52};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd194, 8'd127, 8'd49};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd194, 8'd125, 8'd47};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd180, 8'd111, 8'd36};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd161, 8'd98, 8'd27};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd155, 8'd85, 8'd25};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd163, 8'd69, 8'd18};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd160, 8'd51, 8'd10};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd143, 8'd56, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd143, 8'd115, 8'd94};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd141, 8'd165, 8'd151};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd69, 8'd115, 8'd131};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd65, 8'd111, 8'd126};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd54, 8'd100, 8'd113};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd50, 8'd97, 8'd107};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd51, 8'd98, 8'd108};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd33, 8'd79, 8'd94};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd32, 8'd77, 8'd98};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd45, 8'd90, 8'd113};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd82, 8'd122, 8'd130};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd144, 8'd177, 8'd184};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd158, 8'd182, 8'd194};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd98, 8'd133, 8'd153};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd40, 8'd82, 8'd104};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd41, 8'd88, 8'd108};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd37, 8'd86, 8'd101};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd43, 8'd93, 8'd102};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd45, 8'd94, 8'd109};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd37, 8'd89, 8'd103};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd55, 8'd103, 8'd113};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd100, 8'd134, 8'd136};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd162, 8'd165, 8'd154};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd126, 8'd90, 8'd64};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd133, 8'd58, 8'd18};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd164, 8'd64, 8'd14};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd154, 8'd71, 8'd21};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd158, 8'd88, 8'd28};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd170, 8'd112, 8'd39};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd192, 8'd136, 8'd53};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd216, 8'd155, 8'd66};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd233, 8'd170, 8'd77};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd236, 8'd182, 8'd84};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd233, 8'd190, 8'd88};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd250, 8'd201, 8'd109};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd245, 8'd194, 8'd102};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd227, 8'd185, 8'd99};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd184, 8'd164, 8'd95};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd125, 8'd121, 8'd73};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd98, 8'd91, 8'd45};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd134, 8'd102, 8'd43};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd191, 8'd133, 8'd59};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd190, 8'd119, 8'd39};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd175, 8'd95, 8'd26};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd156, 8'd61, 8'd13};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd126, 8'd31, 8'd1};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd98, 8'd16, 8'd2};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd117, 8'd67, 8'd60};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd164, 8'd146, 8'd142};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd171, 8'd176, 8'd172};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd106, 8'd110, 8'd113};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd97, 8'd86, 8'd80};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd123, 8'd85, 8'd64};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd143, 8'd65, 8'd29};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd171, 8'd57, 8'd7};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd200, 8'd75, 8'd11};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd196, 8'd83, 8'd3};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd204, 8'd106, 8'd17};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd229, 8'd122, 8'd18};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd235, 8'd131, 8'd20};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd243, 8'd140, 8'd19};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd245, 8'd146, 8'd16};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd245, 8'd149, 8'd11};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd245, 8'd152, 8'd12};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd250, 8'd159, 8'd19};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd254, 8'd163, 8'd23};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd247, 8'd170, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd247, 8'd172, 8'd29};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd244, 8'd172, 8'd28};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd237, 8'd170, 8'd27};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd234, 8'd171, 8'd32};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd240, 8'd180, 8'd47};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd254, 8'd196, 8'd70};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd86};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd254, 8'd179, 8'd77};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd242, 8'd158, 8'd62};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd196, 8'd98, 8'd9};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd206, 8'd97, 8'd15};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd227, 8'd112, 8'd31};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd219, 8'd104, 8'd21};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd228, 8'd117, 8'd28};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd219, 8'd111, 8'd20};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd224, 8'd114, 8'd17};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd222, 8'd112, 8'd14};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd218, 8'd111, 8'd7};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd219, 8'd115, 8'd4};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd224, 8'd123, 8'd5};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd235, 8'd137, 8'd12};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd247, 8'd150, 8'd20};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd253, 8'd159, 8'd27};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd40};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd36};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd31};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd251, 8'd163, 8'd27};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd247, 8'd166, 8'd25};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd247, 8'd171, 8'd26};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd176, 8'd27};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd251, 8'd180, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd27};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd26};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd251, 8'd186, 8'd22};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd240, 8'd184, 8'd25};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd230, 8'd184, 8'd47};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd228, 8'd193, 8'd91};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd236, 8'd208, 8'd143};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd245, 8'd222, 8'd180};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd63: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd187};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd251, 8'd211, 8'd160};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd245, 8'd166, 8'd63};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd245, 8'd167, 8'd56};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd245, 8'd172, 8'd44};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd247, 8'd181, 8'd35};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd251, 8'd188, 8'd31};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd250, 8'd191, 8'd25};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd244, 8'd187, 8'd18};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd237, 8'd183, 8'd13};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd47};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd38};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd27};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd254, 8'd160, 8'd26};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd32};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd34};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd34};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd243, 8'd126, 8'd21};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd237, 8'd120, 8'd17};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd229, 8'd109, 8'd12};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd224, 8'd103, 8'd10};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd222, 8'd98, 8'd12};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd217, 8'd90, 8'd9};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd211, 8'd81, 8'd5};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd204, 8'd74, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd220, 8'd95, 8'd5};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd198, 8'd85, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd218, 8'd129, 8'd29};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd249, 8'd182, 8'd75};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd239, 8'd192, 8'd74};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd236, 8'd200, 8'd77};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd251, 8'd222, 8'd92};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd254, 8'd227, 8'd94};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd64};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd48};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd244, 8'd183, 8'd32};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd237, 8'd179, 8'd20};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd239, 8'd175, 8'd17};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd244, 8'd164, 8'd13};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd245, 8'd148, 8'd5};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd242, 8'd135, 8'd0};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd255, 8'd133, 8'd16};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd255, 8'd130, 8'd17};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd245, 8'd124, 8'd20};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd228, 8'd113, 8'd22};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd210, 8'd99, 8'd20};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd191, 8'd82, 8'd17};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd176, 8'd67, 8'd11};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd166, 8'd58, 8'd9};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd156, 8'd24, 8'd0};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd142, 8'd51, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd113, 8'd79, 8'd67};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd94, 8'd94, 8'd94};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd118, 8'd121, 8'd128};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd182, 8'd167, 8'd172};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd177, 8'd144, 8'd139};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd92, 8'd46, 8'd31};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd101, 8'd23, 8'd11};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd132, 8'd39, 8'd6};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd166, 8'd65, 8'd9};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd176, 8'd86, 8'd23};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd161, 8'd97, 8'd36};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd155, 8'd103, 8'd43};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd178, 8'd120, 8'd47};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd211, 8'd139, 8'd54};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd221, 8'd157, 8'd67};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd223, 8'd166, 8'd79};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd229, 8'd178, 8'd97};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd230, 8'd187, 8'd109};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd229, 8'd190, 8'd113};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd223, 8'd185, 8'd104};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd217, 8'd177, 8'd90};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd212, 8'd171, 8'd81};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd204, 8'd150, 8'd54};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd179, 8'd131, 8'd46};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd158, 8'd98, 8'd28};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd167, 8'd73, 8'd19};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd158, 8'd39, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd156, 8'd53, 8'd20};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd135, 8'd91, 8'd62};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd147, 8'd160, 8'd132};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd87, 8'd132, 8'd151};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd85, 8'd131, 8'd146};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd70, 8'd116, 8'd129};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd57, 8'd104, 8'd114};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd59, 8'd105, 8'd118};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd42, 8'd88, 8'd104};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd44, 8'd89, 8'd110};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd51, 8'd95, 8'd120};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd75, 8'd119, 8'd128};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd114, 8'd148, 8'd157};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd205, 8'd224, 8'd230};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd220, 8'd225, 8'd228};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd97, 8'd126, 8'd140};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd75, 8'd113, 8'd134};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd50, 8'd95, 8'd118};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd38, 8'd85, 8'd105};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd46, 8'd94, 8'd106};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd54, 8'd101, 8'd107};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd40, 8'd98, 8'd120};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd55, 8'd111, 8'd128};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd76, 8'd123, 8'd131};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd101, 8'd127, 8'd124};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd159, 8'd153, 8'd137};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd117, 8'd72, 8'd41};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd142, 8'd61, 8'd18};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd163, 8'd61, 8'd12};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd176, 8'd77, 8'd46};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd176, 8'd97, 8'd54};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd184, 8'd130, 8'd68};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd201, 8'd162, 8'd85};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd225, 8'd188, 8'd100};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd243, 8'd206, 8'd115};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd249, 8'd221, 8'd122};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd248, 8'd229, 8'd127};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd137};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd113};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd112};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd132};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd216, 8'd186, 8'd122};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd165, 8'd136, 8'd76};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd166, 8'd118, 8'd42};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd201, 8'd132, 8'd37};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd187, 8'd121, 8'd25};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd178, 8'd99, 8'd22};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd148, 8'd53, 8'd5};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd121, 8'd22, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd104, 8'd24, 8'd17};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd150, 8'd100, 8'd99};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd191, 8'd180, 8'd174};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd148, 8'd161, 8'd151};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd102, 8'd100, 8'd101};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd122, 8'd105, 8'd95};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd119, 8'd72, 8'd46};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd133, 8'd45, 8'd5};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd179, 8'd60, 8'd4};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd204, 8'd77, 8'd8};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd205, 8'd95, 8'd10};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd205, 8'd115, 8'd19};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd235, 8'd131, 8'd18};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd239, 8'd139, 8'd19};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd245, 8'd146, 8'd17};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd246, 8'd153, 8'd14};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd246, 8'd155, 8'd12};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd249, 8'd160, 8'd16};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd27};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd35};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd249, 8'd176, 8'd37};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd253, 8'd182, 8'd42};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd53};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd65};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd75};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd72};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd240, 8'd189, 8'd62};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd225, 8'd175, 8'd52};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd248, 8'd165, 8'd61};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd225, 8'd132, 8'd36};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd175, 8'd67, 8'd0};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd192, 8'd71, 8'd0};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd210, 8'd80, 8'd4};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd192, 8'd61, 8'd0};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd209, 8'd80, 8'd0};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd214, 8'd88, 8'd3};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd213, 8'd94, 8'd0};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd221, 8'd103, 8'd5};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd234, 8'd118, 8'd15};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd247, 8'd135, 8'd25};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd31};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd32};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd28};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd237, 8'd168, 8'd29};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd239, 8'd170, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd244, 8'd176, 8'd33};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd249, 8'd178, 8'd34};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd250, 8'd180, 8'd33};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd250, 8'd180, 8'd32};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd248, 8'd178, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd247, 8'd176, 8'd26};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd0};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd254, 8'd165, 8'd19};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd254, 8'd175, 8'd57};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd111};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd168};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd218};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd64: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd242, 8'd232, 8'd183};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd226, 8'd195, 8'd112};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd240, 8'd204, 8'd108};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd157};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd192};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd180};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd252, 8'd225, 8'd158};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd239, 8'd204, 8'd120};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd229, 8'd187, 8'd79};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd230, 8'd177, 8'd47};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd238, 8'd177, 8'd24};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd252, 8'd184, 8'd13};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd9};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd25};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd25};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd253, 8'd171, 8'd27};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd249, 8'd170, 8'd25};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd244, 8'd169, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd237, 8'd166, 8'd22};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd232, 8'd164, 8'd21};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd229, 8'd162, 8'd19};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd19};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd131, 8'd14};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd245, 8'd121, 8'd9};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd234, 8'd111, 8'd8};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd224, 8'd103, 8'd10};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd214, 8'd96, 8'd9};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd201, 8'd84, 8'd5};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd192, 8'd76, 8'd1};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd210, 8'd84, 8'd10};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd188, 8'd68, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd184, 8'd77, 8'd0};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd246, 8'd155, 8'd64};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd243, 8'd169, 8'd60};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd236, 8'd182, 8'd50};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd245, 8'd204, 8'd52};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd244, 8'd211, 8'd46};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd59};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd251, 8'd221, 8'd65};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd72};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd74};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd67};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd252, 8'd190, 8'd55};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd252, 8'd175, 8'd43};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd252, 8'd169, 8'd39};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd237, 8'd144, 8'd15};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd238, 8'd141, 8'd11};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd239, 8'd137, 8'd9};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd236, 8'd132, 8'd11};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd227, 8'd122, 8'd13};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd205, 8'd104, 8'd14};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd180, 8'd82, 8'd11};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd160, 8'd66, 8'd5};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd148, 8'd50, 8'd3};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd144, 8'd41, 8'd10};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd134, 8'd47, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd137, 8'd99, 8'd88};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd98, 8'd114, 8'd101};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd134, 8'd167, 8'd156};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd172, 8'd176, 8'd177};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd143, 8'd110, 8'd121};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd113, 8'd12, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd130, 8'd21, 8'd0};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd157, 8'd48, 8'd15};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd182, 8'd85, 8'd32};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd193, 8'd111, 8'd37};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd197, 8'd122, 8'd29};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd211, 8'd129, 8'd27};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd227, 8'd136, 8'd31};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd228, 8'd171, 8'd56};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd236, 8'd183, 8'd81};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd245, 8'd198, 8'd116};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd251, 8'd212, 8'd147};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd248, 8'd218, 8'd156};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd238, 8'd214, 8'd144};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd223, 8'd205, 8'd121};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd214, 8'd198, 8'd103};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd206, 8'd177, 8'd107};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd184, 8'd148, 8'd86};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd174, 8'd121, 8'd69};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd163, 8'd87, 8'd38};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd160, 8'd74, 8'd27};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd144, 8'd69, 8'd29};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd126, 8'd80, 8'd54};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd160, 8'd138, 8'd124};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd121, 8'd156, 8'd178};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd76, 8'd122, 8'd138};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd59, 8'd116, 8'd127};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd53, 8'd105, 8'd118};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd60, 8'd99, 8'd116};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd67, 8'd99, 8'd120};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd50, 8'd88, 8'd109};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd51, 8'd98, 8'd118};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd79, 8'd112, 8'd129};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd120, 8'd148, 8'd162};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd180, 8'd200, 8'd209};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd156, 8'd182, 8'd199};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd101, 8'd140, 8'd171};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd80, 8'd120, 8'd155};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd45, 8'd81, 8'd105};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd61, 8'd94, 8'd109};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd55, 8'd98, 8'd107};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd63, 8'd113, 8'd122};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd54, 8'd108, 8'd136};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd66, 8'd124, 8'd146};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd77, 8'd134, 8'd145};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd123, 8'd153, 8'd155};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd159, 8'd146, 8'd137};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd114, 8'd59, 8'd38};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd140, 8'd58, 8'd21};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd157, 8'd66, 8'd19};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd163, 8'd85, 8'd36};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd182, 8'd109, 8'd56};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd209, 8'd145, 8'd84};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd231, 8'd178, 8'd112};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd243, 8'd200, 8'd131};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd248, 8'd215, 8'd144};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd249, 8'd225, 8'd155};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd250, 8'd230, 8'd161};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd247, 8'd248, 8'd146};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd134};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd254, 8'd212, 8'd104};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd245, 8'd179, 8'd69};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd238, 8'd160, 8'd51};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd238, 8'd160, 8'd51};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd234, 8'd166, 8'd57};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd229, 8'd167, 8'd58};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd230, 8'd121, 8'd28};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd174, 8'd61, 8'd0};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd143, 8'd37, 8'd0};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd116, 8'd38, 8'd26};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd94, 8'd56, 8'd55};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd127, 8'd123, 8'd122};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd148, 8'd163, 8'd156};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd110, 8'd130, 8'd119};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd102, 8'd123, 8'd108};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd130, 8'd93, 8'd74};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd161, 8'd60, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd179, 8'd51, 8'd4};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd185, 8'd67, 8'd3};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd193, 8'd91, 8'd7};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd211, 8'd103, 8'd4};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd228, 8'd106, 8'd0};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd230, 8'd133, 8'd0};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd242, 8'd146, 8'd8};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd246, 8'd155, 8'd22};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd241, 8'd158, 8'd26};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd237, 8'd167, 8'd35};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd246, 8'd188, 8'd54};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd71};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd79};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd245, 8'd212, 8'd73};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd77};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd245, 8'd213, 8'd68};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd225, 8'd190, 8'd44};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd234, 8'd191, 8'd53};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd244, 8'd186, 8'd63};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd226, 8'd155, 8'd49};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd231, 8'd151, 8'd54};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd227, 8'd148, 8'd45};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd187, 8'd99, 8'd1};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd179, 8'd75, 8'd0};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd200, 8'd81, 8'd0};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd205, 8'd80, 8'd0};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd206, 8'd84, 8'd1};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd213, 8'd97, 8'd12};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd214, 8'd103, 8'd14};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd234, 8'd123, 8'd8};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd237, 8'd126, 8'd11};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd242, 8'd133, 8'd14};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd246, 8'd142, 8'd19};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd252, 8'd150, 8'd22};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd28};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd31};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd32};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd241, 8'd176, 8'd58};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd241, 8'd180, 8'd38};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd244, 8'd186, 8'd14};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd244, 8'd190, 8'd0};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd245, 8'd188, 8'd0};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd243, 8'd182, 8'd13};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd241, 8'd174, 8'd41};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd61};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd233, 8'd191, 8'd93};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd239, 8'd206, 8'd125};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd247, 8'd230, 8'd178};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd254, 8'd248, 8'd224};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd249, 8'd255, 8'd224};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd241, 8'd243, 8'd178};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd250, 8'd238, 8'd152};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd251, 8'd220, 8'd127};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd224, 8'd181, 8'd89};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd65: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd244, 8'd238, 8'd186};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd228, 8'd198, 8'd112};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd220, 8'd178, 8'd70};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd231, 8'd194, 8'd87};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd243, 8'd218, 8'd118};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd243, 8'd218, 8'd138};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd251, 8'd229, 8'd156};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd252, 8'd245, 8'd226};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd191};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd149};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd249, 8'd195, 8'd105};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd242, 8'd175, 8'd70};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd49};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd252, 8'd176, 8'd12};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd15};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd19};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd23};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd23};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd20};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd17};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd228, 8'd157, 8'd41};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd225, 8'd150, 8'd35};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd223, 8'd139, 8'd27};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd225, 8'd130, 8'd22};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd230, 8'd123, 8'd19};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd232, 8'd114, 8'd14};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd230, 8'd103, 8'd6};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd227, 8'd94, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd214, 8'd89, 8'd9};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd204, 8'd85, 8'd5};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd192, 8'd83, 8'd1};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd232, 8'd136, 8'd49};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd248, 8'd169, 8'd66};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd234, 8'd172, 8'd49};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd230, 8'd181, 8'd40};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd235, 8'd191, 8'd40};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd245, 8'd203, 8'd55};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd249, 8'd209, 8'd62};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd70};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd77};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd77};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd78};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd79};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd80};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd57};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd249, 8'd165, 8'd33};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd238, 8'd149, 8'd21};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd223, 8'd132, 8'd17};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd204, 8'd112, 8'd13};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd181, 8'd90, 8'd7};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd164, 8'd76, 8'd4};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd152, 8'd61, 8'd4};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd143, 8'd44, 8'd2};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd135, 8'd44, 8'd23};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd131, 8'd83, 8'd69};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd96, 8'd99, 8'd88};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd115, 8'd142, 8'd135};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd170, 8'd178, 8'd181};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd178, 8'd158, 8'd170};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd115, 8'd39, 8'd25};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd118, 8'd30, 8'd8};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd140, 8'd41, 8'd2};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd178, 8'd82, 8'd21};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd211, 8'd126, 8'd43};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd224, 8'd148, 8'd50};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd227, 8'd150, 8'd44};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd230, 8'd145, 8'd39};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd227, 8'd159, 8'd48};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd232, 8'd169, 8'd64};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd240, 8'd185, 8'd92};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd247, 8'd200, 8'd118};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd254, 8'd213, 8'd134};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd254, 8'd219, 8'd137};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd134};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd252, 8'd221, 8'd128};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd230, 8'd194, 8'd118};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd208, 8'd164, 8'd99};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd190, 8'd133, 8'd78};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd167, 8'd91, 8'd41};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd156, 8'd70, 8'd23};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd143, 8'd70, 8'd29};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd142, 8'd96, 8'd70};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd184, 8'd162, 8'd148};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd123, 8'd156, 8'd175};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd85, 8'd131, 8'd146};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd66, 8'd123, 8'd134};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd68, 8'd122, 8'd132};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd68, 8'd110, 8'd126};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd76, 8'd111, 8'd131};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd53, 8'd94, 8'd112};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd57, 8'd106, 8'd123};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd64, 8'd105, 8'd125};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd114, 8'd150, 8'd166};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd148, 8'd175, 8'd186};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd143, 8'd176, 8'd193};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd100, 8'd144, 8'd173};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd72, 8'd117, 8'd148};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd55, 8'd93, 8'd116};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd62, 8'd95, 8'd110};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd68, 8'd108, 8'd118};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd69, 8'd117, 8'd129};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd66, 8'd120, 8'd148};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd67, 8'd125, 8'd145};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd84, 8'd138, 8'd148};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd125, 8'd154, 8'd152};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd161, 8'd147, 8'd134};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd116, 8'd60, 8'd35};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd147, 8'd68, 8'd29};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd159, 8'd71, 8'd21};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd160, 8'd93, 8'd41};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd182, 8'd120, 8'd63};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd218, 8'd161, 8'd94};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd244, 8'd196, 8'd120};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd135};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd141};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd144};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd254, 8'd230, 8'd144};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd234, 8'd201, 8'd98};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd242, 8'd199, 8'd94};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd247, 8'd189, 8'd79};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd247, 8'd174, 8'd61};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd249, 8'd168, 8'd53};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd250, 8'd168, 8'd56};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd243, 8'd165, 8'd57};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd233, 8'd156, 8'd52};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd205, 8'd109, 8'd23};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd150, 8'd51, 8'd0};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd128, 8'd35, 8'd2};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd125, 8'd58, 8'd50};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd107, 8'd78, 8'd80};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd100, 8'd104, 8'd105};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd84, 8'd104, 8'd102};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd44, 8'd67, 8'd59};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd84, 8'd91, 8'd73};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd111, 8'd69, 8'd44};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd149, 8'd50, 8'd11};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd173, 8'd52, 8'd0};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd185, 8'd78, 8'd6};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd199, 8'd110, 8'd18};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd221, 8'd128, 8'd22};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd240, 8'd135, 8'd18};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd240, 8'd158, 8'd22};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd252, 8'd174, 8'd38};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd255, 8'd188, 8'd55};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd61};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd254, 8'd197, 8'd64};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd78};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd85};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd85};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd249, 8'd224, 8'd82};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd236, 8'd207, 8'd69};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd241, 8'd202, 8'd71};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd242, 8'd194, 8'd70};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd237, 8'd177, 8'd63};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd212, 8'd143, 8'd40};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd186, 8'd110, 8'd14};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd198, 8'd117, 8'd26};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd208, 8'd114, 8'd52};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd179, 8'd77, 8'd15};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd180, 8'd64, 8'd3};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd203, 8'd78, 8'd12};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd211, 8'd80, 8'd8};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd214, 8'd87, 8'd6};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd224, 8'd105, 8'd13};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd229, 8'd115, 8'd18};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd227, 8'd128, 8'd37};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd233, 8'd136, 8'd39};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd241, 8'd150, 8'd45};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd248, 8'd163, 8'd46};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd251, 8'd172, 8'd41};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd249, 8'd177, 8'd33};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd245, 8'd176, 8'd23};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd241, 8'd175, 8'd18};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd1};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd3};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd249, 8'd164, 8'd11};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd237, 8'd168, 8'd29};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd233, 8'd178, 8'd61};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd236, 8'd193, 8'd99};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd240, 8'd208, 8'd135};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd245, 8'd216, 8'd156};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd191};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd179};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd244, 8'd215, 8'd155};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd246, 8'd210, 8'd122};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd88};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd240, 8'd197, 8'd58};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd233, 8'd184, 8'd55};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd239, 8'd183, 8'd72};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd66: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd250, 8'd249, 8'd203};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd241, 8'd216, 8'd132};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd215, 8'd168, 8'd52};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd214, 8'd156, 8'd23};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd241, 8'd180, 8'd40};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd109};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd245, 8'd209, 8'd97};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd230, 8'd209, 8'd90};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd230, 8'd221, 8'd102};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd240, 8'd239, 8'd133};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd252, 8'd249, 8'd170};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd196};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd210};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd201};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd253, 8'd222, 8'd178};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd247, 8'd213, 8'd165};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd242, 8'd200, 8'd82};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd242, 8'd193, 8'd75};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd240, 8'd184, 8'd61};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd242, 8'd174, 8'd47};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd247, 8'd169, 8'd35};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd27};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd25};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd24};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd17};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd248, 8'd167, 8'd13};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd241, 8'd155, 8'd10};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd235, 8'd144, 8'd11};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd231, 8'd135, 8'd14};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd227, 8'd125, 8'd15};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd218, 8'd112, 8'd12};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd212, 8'd103, 8'd8};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd203, 8'd81, 8'd0};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd201, 8'd85, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd183, 8'd72, 8'd0};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd196, 8'd97, 8'd12};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd237, 8'd150, 8'd57};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd226, 8'd152, 8'd45};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd220, 8'd155, 8'd35};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd224, 8'd165, 8'd35};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd241, 8'd184, 8'd51};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd253, 8'd200, 8'd68};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd86};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd92};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd254, 8'd220, 8'd87};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd248, 8'd215, 8'd84};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd253, 8'd220, 8'd91};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd100};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd85};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd77};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd66};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd58};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd245, 8'd174, 8'd50};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd226, 8'd150, 8'd38};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd201, 8'd123, 8'd25};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd184, 8'd105, 8'd13};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd163, 8'd84, 8'd9};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd145, 8'd52, 8'd0};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd137, 8'd44, 8'd11};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd135, 8'd74, 8'd56};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd119, 8'd102, 8'd94};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd104, 8'd116, 8'd114};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd135, 8'd146, 8'd152};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd147, 8'd145, 8'd159};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd117, 8'd83, 8'd73};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd116, 8'd59, 8'd39};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd134, 8'd51, 8'd7};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd176, 8'd82, 8'd10};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd217, 8'd130, 8'd33};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd238, 8'd161, 8'd53};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd242, 8'd170, 8'd60};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd243, 8'd169, 8'd62};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd250, 8'd169, 8'd61};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd243, 8'd169, 8'd60};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd237, 8'd171, 8'd61};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd233, 8'd175, 8'd67};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd236, 8'd181, 8'd78};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd244, 8'd192, 8'd93};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd254, 8'd201, 8'd109};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd117};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd243, 8'd192, 8'd109};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd224, 8'd170, 8'd98};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd203, 8'd139, 8'd78};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd174, 8'd97, 8'd43};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd153, 8'd70, 8'd20};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd141, 8'd68, 8'd27};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd148, 8'd101, 8'd75};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd187, 8'd161, 8'd148};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd135, 8'd164, 8'd180};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd103, 8'd145, 8'd157};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd77, 8'd134, 8'd143};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd79, 8'd136, 8'd145};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd81, 8'd127, 8'd142};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd87, 8'd125, 8'd144};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd61, 8'd104, 8'd121};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd61, 8'd113, 8'd127};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd54, 8'd104, 8'd129};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd106, 8'd151, 8'd172};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd117, 8'd150, 8'd165};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd200, 8'd231, 8'd234};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd124, 8'd166, 8'd180};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd91, 8'd143, 8'd167};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd63, 8'd113, 8'd140};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd65, 8'd106, 8'd126};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd65, 8'd101, 8'd113};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd81, 8'd119, 8'd130};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd76, 8'd122, 8'd137};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd74, 8'd128, 8'd154};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd71, 8'd128, 8'd145};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd97, 8'd148, 8'd152};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd140, 8'd163, 8'd157};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd159, 8'd140, 8'd125};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd119, 8'd62, 8'd33};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd150, 8'd73, 8'd29};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd160, 8'd77, 8'd23};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd163, 8'd106, 8'd51};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd185, 8'd129, 8'd68};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd214, 8'd162, 8'd89};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd238, 8'd188, 8'd103};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd246, 8'd200, 8'd104};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd244, 8'd201, 8'd97};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd239, 8'd198, 8'd92};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd236, 8'd195, 8'd89};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd244, 8'd170, 8'd65};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd249, 8'd176, 8'd65};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd253, 8'd181, 8'd63};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd59};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd61};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd60};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd243, 8'd155, 8'd49};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd224, 8'd132, 8'd33};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd180, 8'd99, 8'd20};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd145, 8'd60, 8'd3};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd129, 8'd50, 8'd19};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd128, 8'd74, 8'd64};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd117, 8'd97, 8'd96};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd103, 8'd109, 8'd109};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd85, 8'd101, 8'd98};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd63, 8'd80, 8'd74};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd94, 8'd80, 8'd53};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd122, 8'd70, 8'd31};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd157, 8'd66, 8'd11};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd186, 8'd82, 8'd11};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd203, 8'd115, 8'd28};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd219, 8'd150, 8'd47};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd243, 8'd174, 8'd57};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd57};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd67};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd80};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd86};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd86};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd254, 8'd215, 8'd84};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd88};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd249, 8'd218, 8'd91};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd243, 8'd214, 8'd86};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd244, 8'd226, 8'd82};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd82};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd241, 8'd193, 8'd83};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd213, 8'd146, 8'd57};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd199, 8'd117, 8'd41};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd209, 8'd123, 8'd48};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd198, 8'd112, 8'd35};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd183, 8'd100, 8'd20};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd181, 8'd75, 8'd33};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd172, 8'd61, 8'd15};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd188, 8'd69, 8'd11};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd214, 8'd91, 8'd21};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd222, 8'd98, 8'd10};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd221, 8'd102, 8'd0};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd227, 8'd116, 8'd0};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd232, 8'd127, 8'd0};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd248, 8'd141, 8'd11};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd249, 8'd145, 8'd14};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd250, 8'd152, 8'd15};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd252, 8'd161, 8'd20};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd253, 8'd168, 8'd23};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd252, 8'd174, 8'd22};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd251, 8'd178, 8'd23};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd249, 8'd180, 8'd24};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd254, 8'd171, 8'd15};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd253, 8'd177, 8'd42};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd254, 8'd185, 8'd90};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd144};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd189};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd254, 8'd246, 8'd183};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd240, 8'd233, 8'd155};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd230, 8'd222, 8'd137};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd215, 8'd203, 8'd81};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd240, 8'd207, 8'd102};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd100};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd72};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd31};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd230, 8'd169, 8'd0};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd214, 8'd163, 8'd22};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd247, 8'd204, 8'd100};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd67: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd181};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd241, 8'd192, 8'd90};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd229, 8'd155, 8'd20};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd250, 8'd161, 8'd7};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd237, 8'd180, 8'd77};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd244, 8'd196, 8'd86};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd248, 8'd213, 8'd93};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd240, 8'd217, 8'd89};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd229, 8'd209, 8'd84};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd231, 8'd205, 8'd92};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd249, 8'd213, 8'd116};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd136};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd254, 8'd228, 8'd151};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd253, 8'd231, 8'd156};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd251, 8'd236, 8'd169};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd251, 8'd242, 8'd183};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd250, 8'd250, 8'd200};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd249, 8'd255, 8'd214};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd248, 8'd255, 8'd226};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd248, 8'd255, 8'd230};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd222};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd254, 8'd239, 8'd206};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd245, 8'd225, 8'd175};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd236, 8'd209, 8'd140};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd230, 8'd196, 8'd106};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd227, 8'd189, 8'd78};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd230, 8'd186, 8'd61};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd232, 8'd186, 8'd51};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd253, 8'd161, 8'd0};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd247, 8'd155, 8'd0};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd240, 8'd147, 8'd0};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd237, 8'd142, 8'd0};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd237, 8'd140, 8'd7};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd232, 8'd137, 8'd11};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd225, 8'd129, 8'd9};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd219, 8'd122, 8'd7};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd220, 8'd107, 8'd15};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd205, 8'd95, 8'd8};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd186, 8'd79, 8'd0};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd175, 8'd75, 8'd0};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd210, 8'd119, 8'd38};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd210, 8'd126, 8'd38};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd210, 8'd134, 8'd36};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd205, 8'd132, 8'd27};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd226, 8'd153, 8'd42};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd239, 8'd172, 8'd59};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd80};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd94};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd99};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd242, 8'd221, 8'd94};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd232, 8'd217, 8'd92};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd226, 8'd215, 8'd91};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd245, 8'd222, 8'd84};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd248, 8'd221, 8'd82};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd80};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd79};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd77};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd245, 8'd186, 8'd66};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd225, 8'd161, 8'd51};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd212, 8'd145, 8'd40};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd179, 8'd109, 8'd21};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd159, 8'd76, 8'd6};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd154, 8'd63, 8'd18};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd139, 8'd67, 8'd43};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd131, 8'd94, 8'd85};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd88, 8'd84, 8'd83};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd86, 8'd97, 8'd103};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd88, 8'd100, 8'd112};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd97};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd113, 8'd83, 8'd59};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd138, 8'd68, 8'd17};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd171, 8'd82, 8'd0};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd199, 8'd111, 8'd5};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd218, 8'd141, 8'd25};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd235, 8'd168, 8'd53};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd251, 8'd184, 8'd77};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd70};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd63};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd250, 8'd176, 8'd51};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd241, 8'd174, 8'd44};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd237, 8'd172, 8'd46};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd237, 8'd170, 8'd57};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd71};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd244, 8'd168, 8'd80};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd233, 8'd168, 8'd76};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd219, 8'd154, 8'd74};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd201, 8'd132, 8'd65};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd181, 8'd102, 8'd45};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd160, 8'd74, 8'd23};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd140, 8'd65, 8'd23};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd139, 8'd85, 8'd57};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd154, 8'd121, 8'd104};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd158, 8'd180, 8'd191};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd126, 8'd163, 8'd171};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd93, 8'd146, 8'd152};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd77, 8'd134, 8'd143};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd95, 8'd143, 8'd157};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd92, 8'd134, 8'd150};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd72, 8'd118, 8'd133};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd60, 8'd112, 8'd123};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd54, 8'd114, 8'd142};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd92, 8'd144, 8'd168};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd104, 8'd146, 8'd162};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd190, 8'd219, 8'd227};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd157, 8'd171, 8'd172};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd157, 8'd179, 8'd177};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd162, 8'd188, 8'd185};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd182, 8'd200, 8'd200};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd224, 8'd225, 8'd230};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd166, 8'd204, 8'd207};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd107, 8'd155, 8'd169};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd75, 8'd131, 8'd154};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd59, 8'd113, 8'd137};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd68, 8'd111, 8'd127};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd75, 8'd111, 8'd123};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd89, 8'd127, 8'd140};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd83, 8'd126, 8'd143};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd72, 8'd124, 8'd148};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd83, 8'd136, 8'd150};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd117, 8'd158, 8'd160};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd164, 8'd176, 8'd166};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd148, 8'd120, 8'd99};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd123, 8'd60, 8'd27};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd144, 8'd66, 8'd18};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd158, 8'd77, 8'd21};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd169, 8'd106, 8'd52};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd183, 8'd122, 8'd59};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd205, 8'd143, 8'd66};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd221, 8'd160, 8'd69};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd230, 8'd167, 8'd62};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd232, 8'd169, 8'd55};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd235, 8'd170, 8'd50};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd236, 8'd172, 8'd49};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd58};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd57};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd54};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd250, 8'd186, 8'd52};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd250, 8'd188, 8'd55};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd243, 8'd173, 8'd51};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd220, 8'd138, 8'd28};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd196, 8'd104, 8'd5};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd152, 8'd74, 8'd0};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd146, 8'd66, 8'd5};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd129, 8'd55, 8'd18};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd107, 8'd55, 8'd34};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd96, 8'd72, 8'd60};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd97, 8'd93, 8'd81};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd104, 8'd105, 8'd91};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd110, 8'd107, 8'd92};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd122, 8'd86, 8'd50};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd147, 8'd87, 8'd37};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd179, 8'd96, 8'd26};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd203, 8'd119, 8'd33};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd220, 8'd150, 8'd54};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd233, 8'd181, 8'd71};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd249, 8'd204, 8'd79};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd80};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd96};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd99};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd254, 8'd225, 8'd97};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd245, 8'd218, 8'd89};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd240, 8'd215, 8'd88};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd244, 8'd219, 8'd93};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd247, 8'd218, 8'd98};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd244, 8'd213, 8'd97};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd238, 8'd214, 8'd80};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd234, 8'd193, 8'd79};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd221, 8'd157, 8'd70};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd169, 8'd83, 8'd24};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd156, 8'd58, 8'd11};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd199, 8'd101, 8'd52};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd202, 8'd112, 8'd52};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd168, 8'd85, 8'd15};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd155, 8'd56, 8'd0};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd178, 8'd76, 8'd0};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd205, 8'd101, 8'd4};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd216, 8'd115, 8'd1};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd219, 8'd124, 8'd0};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd232, 8'd142, 8'd4};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd244, 8'd159, 8'd16};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd242, 8'd156, 8'd0};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd240, 8'd157, 8'd0};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd240, 8'd162, 8'd14};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd239, 8'd167, 8'd31};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd239, 8'd173, 8'd51};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd241, 8'd180, 8'd73};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd241, 8'd186, 8'd86};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd242, 8'd189, 8'd95};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd238, 8'd230, 8'd147};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd245, 8'd236, 8'd171};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd207};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd247, 8'd212};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd242, 8'd244, 8'd195};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd194};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd177};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd245, 8'd214, 8'd149};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd241, 8'd204, 8'd124};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd240, 8'd204, 8'd108};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd243, 8'd209, 8'd101};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd246, 8'd215, 8'd98};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd246, 8'd217, 8'd97};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd239, 8'd232, 8'd99};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd251, 8'd217, 8'd107};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd89};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd44};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd238, 8'd159, 8'd0};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd206, 8'd150, 8'd0};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd213, 8'd181, 8'd78};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd251, 8'd237, 8'd188};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd68: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd227};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd160};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd249, 8'd177, 8'd67};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd246, 8'd153, 8'd14};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd228, 8'd134, 8'd20};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd242, 8'd156, 8'd47};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd84};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd112};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd122};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd253, 8'd213, 8'd115};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd244, 8'd209, 8'd105};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd241, 8'd209, 8'd98};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd250, 8'd206, 8'd75};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd249, 8'd210, 8'd83};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd247, 8'd214, 8'd98};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd244, 8'd221, 8'd117};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd240, 8'd227, 8'd135};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd234, 8'd231, 8'd152};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd230, 8'd233, 8'd162};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd226, 8'd235, 8'd170};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd252, 8'd238, 8'd225};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd223};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd218};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd205};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd188};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd251, 8'd243, 8'd170};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd243, 8'd235, 8'd150};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd238, 8'd231, 8'd141};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd249, 8'd209, 8'd121};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd244, 8'd199, 8'd106};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd238, 8'd184, 8'd84};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd236, 8'd170, 8'd60};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd236, 8'd157, 8'd38};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd233, 8'd144, 8'd14};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd227, 8'd129, 8'd0};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd221, 8'd118, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd218, 8'd119, 8'd26};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd185, 8'd86, 8'd1};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd175, 8'd77, 8'd2};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd155, 8'd60, 8'd0};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd171, 8'd79, 8'd12};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd186, 8'd98, 8'd27};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd203, 8'd120, 8'd42};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd189, 8'd107, 8'd25};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd198, 8'd112, 8'd25};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd205, 8'd124, 8'd32};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd223, 8'd151, 8'd49};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd243, 8'd186, 8'd73};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd96};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd109};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd245, 8'd226, 8'd106};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd231, 8'd219, 8'd99};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd241, 8'd222, 8'd93};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd239, 8'd219, 8'd88};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd238, 8'd214, 8'd82};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd240, 8'd211, 8'd81};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd243, 8'd205, 8'd80};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd240, 8'd195, 8'd76};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd233, 8'd181, 8'd69};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd227, 8'd171, 8'd62};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd194, 8'd129, 8'd37};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd185, 8'd109, 8'd33};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd174, 8'd91, 8'd37};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd135, 8'd60, 8'd28};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd118, 8'd69, 8'd52};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd83, 8'd64, 8'd58};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd78, 8'd82, 8'd83};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd85, 8'd98, 8'd104};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd83, 8'd96, 8'd86};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd102, 8'd82, 8'd57};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd138, 8'd77, 8'd23};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd175, 8'd89, 8'd6};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd198, 8'd112, 8'd3};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd212, 8'd138, 8'd17};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd231, 8'd166, 8'd46};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd249, 8'd187, 8'd74};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd65};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd62};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd58};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd55};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd56};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd253, 8'd181, 8'd60};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd246, 8'd167, 8'd64};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd243, 8'd158, 8'd67};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd228, 8'd152, 8'd54};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd211, 8'd139, 8'd54};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd192, 8'd120, 8'd48};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd181, 8'd101, 8'd40};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd163, 8'd78, 8'd23};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd144, 8'd66, 8'd18};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd133, 8'd73, 8'd39};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd125, 8'd80, 8'd57};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd178, 8'd189, 8'd195};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd151, 8'd180, 8'd184};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd113, 8'd160, 8'd166};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd71, 8'd125, 8'd135};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd105, 8'd152, 8'd168};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd97, 8'd139, 8'd155};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd88, 8'd134, 8'd147};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd62, 8'd112, 8'd121};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd57, 8'd120, 8'd151};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd70, 8'd126, 8'd151};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd106, 8'd149, 8'd166};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd151, 8'd181, 8'd191};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd202, 8'd212, 8'd211};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd178, 8'd182, 8'd181};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd204, 8'd200, 8'd199};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd208, 8'd199, 8'd202};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd146, 8'd164, 8'd166};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd147, 8'd173, 8'd172};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd139, 8'd169, 8'd167};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd135, 8'd156, 8'd157};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd153, 8'd160, 8'd166};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd194, 8'd193, 8'd201};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd137, 8'd174, 8'd180};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd100, 8'd148, 8'd162};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd61, 8'd118, 8'd138};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd64, 8'd119, 8'd139};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd69, 8'd113, 8'd126};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd89, 8'd126, 8'd135};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd94, 8'd132, 8'd145};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd89, 8'd132, 8'd151};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd68, 8'd116, 8'd138};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd105, 8'd151, 8'd164};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd140, 8'd170, 8'd170};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd183, 8'd181, 8'd168};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd133, 8'd91, 8'd66};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd128, 8'd56, 8'd18};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd134, 8'd52, 8'd2};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd154, 8'd74, 8'd15};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd168, 8'd91, 8'd35};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd186, 8'd108, 8'd44};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd208, 8'd131, 8'd53};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd230, 8'd151, 8'd58};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd244, 8'd163, 8'd55};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd251, 8'd170, 8'd52};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd51};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd52};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd55};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd254, 8'd179, 8'd54};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd243, 8'd184, 8'd48};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd235, 8'd186, 8'd45};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd234, 8'd187, 8'd49};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd229, 8'd174, 8'd47};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd211, 8'd141, 8'd29};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd187, 8'd108, 8'd5};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd169, 8'd88, 8'd9};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd164, 8'd81, 8'd15};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd142, 8'd61, 8'd14};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd114, 8'd51, 8'd18};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd95, 8'd58, 8'd29};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd91, 8'd65, 8'd38};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd100, 8'd73, 8'd44};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd120, 8'd85, 8'd57};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd137, 8'd79, 8'd39};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd156, 8'd91, 8'd33};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd181, 8'd113, 8'd32};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd205, 8'd139, 8'd43};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd220, 8'd165, 8'd64};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd231, 8'd189, 8'd79};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd242, 8'd207, 8'd87};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd248, 8'd218, 8'd86};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd106};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd249, 8'd224, 8'd106};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd246, 8'd224, 8'd102};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd240, 8'd219, 8'd94};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd243, 8'd217, 8'd94};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd253, 8'd220, 8'd104};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd107};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd254, 8'd205, 8'd103};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd232, 8'd180, 8'd70};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd191, 8'd126, 8'd34};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd174, 8'd93, 8'd27};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd161, 8'd64, 8'd21};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd153, 8'd50, 8'd17};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd162, 8'd62, 8'd26};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd156, 8'd64, 8'd15};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd145, 8'd61, 8'd1};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd148, 8'd63, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd158, 8'd74, 8'd1};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd173, 8'd88, 8'd5};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd185, 8'd105, 8'd10};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd194, 8'd117, 8'd13};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd197, 8'd126, 8'd18};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd209, 8'd143, 8'd33};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd226, 8'd162, 8'd52};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd201, 8'd169, 8'd56};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd209, 8'd181, 8'd72};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd223, 8'd199, 8'd101};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd237, 8'd219, 8'd135};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd249, 8'd236, 8'd168};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd254, 8'd247, 8'd193};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd254, 8'd211};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd218};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd239, 8'd248, 8'd205};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd241, 8'd247, 8'd203};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd243, 8'd245, 8'd195};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd247, 8'd242, 8'd186};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd246, 8'd236, 8'd167};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd244, 8'd228, 8'd150};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd241, 8'd221, 8'd132};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd240, 8'd217, 8'd123};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd244, 8'd205, 8'd104};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd251, 8'd210, 8'd105};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd108};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd107};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd106};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd103};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd250, 8'd214, 8'd102};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd102};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd109};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd248, 8'd190, 8'd83};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd242, 8'd154, 8'd54};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd234, 8'd135, 8'd16};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd223, 8'd135, 8'd1};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd231, 8'd174, 8'd59};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd251, 8'd224, 8'd169};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd69: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd216};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd253, 8'd203, 8'd130};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd233, 8'd160, 8'd55};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd0};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd250, 8'd127, 8'd0};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd238, 8'd125, 8'd21};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd251, 8'd152, 8'd71};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd127};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd159};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd157};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd237, 8'd232, 8'd141};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd114};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd114};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd247, 8'd218, 8'd114};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd113};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd249, 8'd214, 8'd112};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd248, 8'd210, 8'd109};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd247, 8'd208, 8'd107};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd248, 8'd206, 8'd106};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd236, 8'd199, 8'd110};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd242, 8'd206, 8'd120};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd134};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd152};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd165};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd176};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd180};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd182};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd192};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd179};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd161};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd247, 8'd215, 8'd140};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd243, 8'd205, 8'd124};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd236, 8'd192, 8'd103};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd227, 8'd178, 8'd85};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd219, 8'd169, 8'd72};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd228, 8'd146, 8'd60};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd190, 8'd107, 8'd29};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd183, 8'd98, 8'd31};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd163, 8'd77, 8'd18};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd152, 8'd65, 8'd11};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd168, 8'd81, 8'd27};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd182, 8'd96, 8'd35};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd170, 8'd85, 8'd20};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd170, 8'd77, 8'd10};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd189, 8'd99, 8'd23};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd214, 8'd130, 8'd42};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd230, 8'd157, 8'd54};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd66};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd245, 8'd196, 8'd78};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd99};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd113};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd108};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd108};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd106};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd106};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd251, 8'd219, 8'd106};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd246, 8'd208, 8'd99};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd191, 8'd86};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd227, 8'd180, 8'd76};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd211, 8'd145, 8'd61};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd193, 8'd125, 8'd50};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd173, 8'd103, 8'd43};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd135, 8'd68, 8'd26};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd126, 8'd72, 8'd46};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd118, 8'd86, 8'd71};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd105, 8'd95, 8'd86};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd98, 8'd103, 8'd97};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd84, 8'd89, 8'd69};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd104, 8'd79, 8'd49};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd145, 8'd83, 8'd32};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd194, 8'd111, 8'd33};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd228, 8'd147, 8'd42};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd243, 8'd172, 8'd54};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd251, 8'd187, 8'd64};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd75};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd73};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd254, 8'd192, 8'd69};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd252, 8'd193, 8'd63};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd250, 8'd192, 8'd58};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd250, 8'd187, 8'd56};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd250, 8'd181, 8'd60};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd251, 8'd174, 8'd66};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd252, 8'd170, 8'd71};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd239, 8'd155, 8'd56};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd218, 8'd141, 8'd53};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd191, 8'd117, 8'd44};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd180, 8'd101, 8'd35};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd164, 8'd78, 8'd17};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd151, 8'd66, 8'd12};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd146, 8'd75, 8'd33};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd124, 8'd65, 8'd35};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd173, 8'd171, 8'd174};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd177, 8'd195, 8'd197};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd140, 8'd179, 8'd184};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd84, 8'd134, 8'd145};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd111, 8'd157, 8'd173};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd112, 8'd151, 8'd168};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd109, 8'd151, 8'd163};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd76, 8'd123, 8'd129};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd65, 8'd122, 8'd152};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd61, 8'd112, 8'd139};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd112, 8'd153, 8'd173};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd131, 8'd161, 8'd172};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd157};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd147, 8'd132, 8'd125};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd180, 8'd159, 8'd154};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd167, 8'd143, 8'd141};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd181, 8'd161, 8'd163};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd189, 8'd182, 8'd189};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd160, 8'd175, 8'd182};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd141, 8'd166, 8'd170};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd124, 8'd155, 8'd157};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd123, 8'd147, 8'd151};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd129, 8'd139, 8'd148};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd142, 8'd146, 8'd157};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd168, 8'd178, 8'd187};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd192, 8'd211, 8'd217};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd124, 8'd154, 8'd165};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd103, 8'd144, 8'd162};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd61, 8'd113, 8'd135};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd74, 8'd125, 8'd144};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd80, 8'd122, 8'd134};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd104, 8'd141, 8'd149};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd104, 8'd141, 8'd157};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd95, 8'd140, 8'd163};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd82, 8'd123, 8'd145};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd136, 8'd172, 8'd184};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd163, 8'd179, 8'd178};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd181, 8'd164, 8'd148};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd125, 8'd68, 8'd41};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd134, 8'd52, 8'd12};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd134, 8'd47, 8'd0};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd152, 8'd70, 8'd10};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd174, 8'd85, 8'd25};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd193, 8'd106, 8'd37};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd221, 8'd134, 8'd54};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd243, 8'd159, 8'd63};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd64};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd255, 8'd175, 8'd59};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd54};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd52};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd247, 8'd182, 8'd64};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd248, 8'd190, 8'd65};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd243, 8'd195, 8'd61};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd239, 8'd198, 8'd58};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd242, 8'd199, 8'd61};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd244, 8'd193, 8'd66};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd232, 8'd170, 8'd57};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd216, 8'd147, 8'd43};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd213, 8'd131, 8'd55};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd177, 8'd92, 8'd27};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd143, 8'd62, 8'd9};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd132, 8'd65, 8'd23};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd119, 8'd71, 8'd31};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd103, 8'd61, 8'd23};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd111, 8'd59, 8'd22};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd139, 8'd75, 8'd40};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd147, 8'd78, 8'd37};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd164, 8'd100, 8'd38};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd187, 8'd131, 8'd44};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd210, 8'd160, 8'd61};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd226, 8'd180, 8'd82};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd239, 8'd197, 8'd97};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd245, 8'd211, 8'd103};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd250, 8'd221, 8'd103};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd124};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd122};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd115};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd253, 8'd223, 8'd103};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd253, 8'd214, 8'd97};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd95};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd248, 8'd179, 8'd84};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd235, 8'd157, 8'd72};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd214, 8'd118, 8'd42};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd165, 8'd68, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd152, 8'd52, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd158, 8'd59, 8'd17};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd159, 8'd63, 8'd25};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd18};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd140, 8'd54, 8'd7};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd152, 8'd69, 8'd17};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd138, 8'd54, 8'd10};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd165, 8'd83, 8'd33};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd192, 8'd116, 8'd56};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd217, 8'd149, 8'd78};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd241, 8'd177, 8'd103};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd252, 8'd194, 8'd121};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd135};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd154};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd168};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd170};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd171};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd171};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd253, 8'd239, 8'd168};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd243, 8'd237, 8'd163};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd235, 8'd233, 8'd158};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd229, 8'd230, 8'd154};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd213, 8'd133};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd248, 8'd212, 8'd124};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd246, 8'd213, 8'd108};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd244, 8'd214, 8'd94};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd246, 8'd215, 8'd88};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd248, 8'd217, 8'd90};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd218, 8'd95};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd254, 8'd219, 8'd101};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd110};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd104};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd238, 8'd214, 8'd106};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd243, 8'd221, 8'd120};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd139};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd144};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd254, 8'd216, 8'd131};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd245, 8'd200, 8'd117};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd244, 8'd146, 8'd35};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd235, 8'd131, 8'd16};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd244, 8'd134, 8'd11};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd246, 8'd141, 8'd13};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd244, 8'd157, 8'd41};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd129};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd70: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd191};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd233, 8'd195, 8'd120};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd12};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd253, 8'd150, 8'd11};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd247, 8'd133, 8'd9};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd241, 8'd126, 8'd19};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd237, 8'd136, 8'd44};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd243, 8'd168, 8'd87};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd254, 8'd208, 8'd131};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd163};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd252, 8'd236, 8'd161};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd250, 8'd233, 8'd155};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd249, 8'd227, 8'd144};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd249, 8'd222, 8'd133};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd253, 8'd219, 8'd122};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd116};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd113};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd111};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd254, 8'd214, 8'd82};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd252, 8'd212, 8'd81};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd85};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd243, 8'd203, 8'd89};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd240, 8'd201, 8'd96};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd240, 8'd202, 8'd105};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd243, 8'd203, 8'd115};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd243, 8'd206, 8'd118};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd249, 8'd207, 8'd109};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd245, 8'd205, 8'd110};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd242, 8'd205, 8'd117};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd244, 8'd211, 8'd132};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd249, 8'd219, 8'd149};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd251, 8'd226, 8'd162};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd248, 8'd226, 8'd169};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd245, 8'd224, 8'd171};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd250, 8'd184, 8'd106};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd227, 8'd160, 8'd89};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd212, 8'd142, 8'd82};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd189, 8'd113, 8'd64};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd161, 8'd82, 8'd39};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd161, 8'd78, 8'd34};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd144, 8'd61, 8'd11};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd148, 8'd65, 8'd11};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd154, 8'd58, 8'd8};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd179, 8'd83, 8'd23};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd209, 8'd113, 8'd36};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd221, 8'd130, 8'd37};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd223, 8'd138, 8'd31};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd227, 8'd151, 8'd39};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd244, 8'd177, 8'd64};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd85};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd99};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd104};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd116};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd127};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd134};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd126};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd245, 8'd206, 8'd113};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd193, 8'd101};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd234, 8'd164, 8'd92};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd198, 8'd135, 8'd66};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd170, 8'd112, 8'd49};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd145, 8'd92, 8'd42};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd140, 8'd88, 8'd51};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd148, 8'd106, 8'd81};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd112, 8'd90, 8'd69};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd89, 8'd80, 8'd63};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd100, 8'd85, 8'd56};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd112, 8'd74, 8'd38};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd145, 8'd79, 8'd29};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd193, 8'd113, 8'd42};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd231, 8'd157, 8'd62};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd250, 8'd184, 8'd71};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd71};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd70};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd85};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd251, 8'd207, 8'd82};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd242, 8'd198, 8'd73};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd236, 8'd190, 8'd68};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd236, 8'd184, 8'd66};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd240, 8'd180, 8'd66};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd248, 8'd180, 8'd71};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd253, 8'd180, 8'd75};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd243, 8'd157, 8'd58};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd227, 8'd147, 8'd60};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd199, 8'd125, 8'd52};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd187, 8'd108, 8'd42};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd165, 8'd77, 8'd13};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd154, 8'd64, 8'd4};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd158, 8'd76, 8'd28};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd134, 8'd62, 8'd22};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd147, 8'd133, 8'd133};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd199, 8'd207, 8'd209};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd167, 8'd200, 8'd205};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd117, 8'd161, 8'd174};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd115, 8'd156, 8'd174};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd134, 8'd169, 8'd188};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd130, 8'd166, 8'd180};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd103, 8'd144, 8'd150};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd77, 8'd126, 8'd156};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd76, 8'd120, 8'd145};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd121, 8'd158, 8'd177};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd150, 8'd176, 8'd189};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd194, 8'd186, 8'd183};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd159, 8'd144, 8'd137};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd148, 8'd107, 8'd87};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd133, 8'd88, 8'd69};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd185, 8'd134, 8'd117};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd150, 8'd98, 8'd85};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd133, 8'd90, 8'd83};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd138, 8'd110, 8'd106};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd178, 8'd170, 8'd168};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd180, 8'd193, 8'd202};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd152, 8'd175, 8'd181};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd130, 8'd159, 8'd163};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd128, 8'd153, 8'd158};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd133, 8'd147, 8'd156};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd131, 8'd141, 8'd151};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd145, 8'd152};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd125, 8'd153, 8'd157};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd127, 8'd146, 8'd163};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd112, 8'd144, 8'd165};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd76, 8'd121, 8'd144};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd82, 8'd129, 8'd147};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd102, 8'd142, 8'd152};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd116, 8'd150, 8'd159};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd120, 8'd159, 8'd174};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd102, 8'd148, 8'd172};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd115, 8'd147, 8'd170};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd168, 8'd194, 8'd207};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd183, 8'd188, 8'd184};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd159, 8'd128, 8'd110};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd127, 8'd58, 8'd29};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd9};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd148, 8'd54, 8'd2};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd156, 8'd70, 8'd9};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd184, 8'd97, 8'd26};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd200, 8'd117, 8'd41};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd223, 8'd143, 8'd56};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd240, 8'd164, 8'd66};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd246, 8'd175, 8'd67};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd64};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd244, 8'd179, 8'd61};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd242, 8'd180, 8'd61};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd243, 8'd198, 8'd83};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd251, 8'd206, 8'd87};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd84};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd77};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd73};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd253, 8'd193, 8'd73};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd241, 8'd174, 8'd67};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd227, 8'd158, 8'd55};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd195, 8'd120, 8'd55};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd153, 8'd74, 8'd17};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd126, 8'd49, 8'd3};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd124, 8'd61, 8'd20};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd117, 8'd68, 8'd28};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd108, 8'd60, 8'd22};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd126, 8'd63, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd154, 8'd77, 8'd47};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd169, 8'd94, 8'd54};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd183, 8'd121, 8'd60};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd204, 8'd158, 8'd72};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd226, 8'd186, 8'd90};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd243, 8'd200, 8'd108};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd252, 8'd206, 8'd118};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd121};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd120};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd125};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd118};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd253, 8'd211, 8'd103};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd244, 8'd197, 8'd83};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd241, 8'd181, 8'd71};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd238, 8'd160, 8'd62};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd226, 8'd127, 8'd44};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd210, 8'd99, 8'd27};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd195, 8'd53, 8'd15};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd173, 8'd42, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd159, 8'd47, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd147, 8'd53, 8'd1};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd149, 8'd68, 8'd13};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd152, 8'd75, 8'd21};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd150, 8'd70, 8'd19};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd171, 8'd89, 8'd41};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd203, 8'd109, 8'd81};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd227, 8'd139, 8'd99};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd243, 8'd164, 8'd108};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd252, 8'd184, 8'd113};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd126};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd127};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd248, 8'd199, 8'd122};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd250, 8'd202, 8'd128};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd110};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd253, 8'd191, 8'd106};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd252, 8'd193, 8'd103};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd196, 8'd98};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd250, 8'd201, 8'd96};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd250, 8'd207, 8'd94};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd92};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd93};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd97};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd96};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd95};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd94};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd96};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd251, 8'd215, 8'd101};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd105};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd109};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd122};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd245, 8'd222, 8'd129};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd242, 8'd227, 8'd142};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd250, 8'd234, 8'd157};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd156};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd128};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd240, 8'd163, 8'd81};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd226, 8'd132, 8'd45};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd124, 8'd27};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd138, 8'd15};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd251, 8'd152, 8'd6};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd237, 8'd161, 8'd23};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd239, 8'd185, 8'd87};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd177};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd71: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd247, 8'd235, 8'd175};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd223, 8'd188, 8'd60};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd234, 8'd178, 8'd43};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd245, 8'd158, 8'd17};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd247, 8'd134, 8'd0};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd241, 8'd118, 8'd0};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd235, 8'd120, 8'd11};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd233, 8'd138, 8'd46};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd235, 8'd154, 8'd75};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd145};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd254, 8'd230, 8'd144};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd252, 8'd228, 8'd140};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd249, 8'd228, 8'd137};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd247, 8'd228, 8'd134};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd246, 8'd227, 8'd132};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd244, 8'd228, 8'd130};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd244, 8'd229, 8'd128};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd114};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd111};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd226, 8'd103};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd252, 8'd221, 8'd96};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd251, 8'd216, 8'd86};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd251, 8'd215, 8'd79};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd252, 8'd215, 8'd75};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd73};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd89};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd240, 8'd203, 8'd86};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd234, 8'd191, 8'd79};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd230, 8'd181, 8'd78};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd231, 8'd172, 8'd80};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd227, 8'd162, 8'd78};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd222, 8'd150, 8'd74};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd216, 8'd142, 8'd69};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd194, 8'd140, 8'd66};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd197, 8'd139, 8'd75};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd185, 8'd122, 8'd69};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd173, 8'd104, 8'd62};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd159, 8'd85, 8'd46};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd154, 8'd76, 8'd37};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd122, 8'd41, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd148, 8'd66, 8'd18};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd148, 8'd52, 8'd10};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd157, 8'd60, 8'd7};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd178, 8'd77, 8'd7};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd204, 8'd103, 8'd13};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd226, 8'd127, 8'd23};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd236, 8'd144, 8'd33};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd235, 8'd149, 8'd36};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd230, 8'd148, 8'd36};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd236, 8'd165, 8'd75};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd235, 8'd171, 8'd81};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd236, 8'd182, 8'd92};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd243, 8'd199, 8'd112};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd250, 8'd214, 8'd126};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd135};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd133};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd253, 8'd215, 8'd130};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd254, 8'd180, 8'd117};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd212, 8'd151, 8'd88};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd180, 8'd130, 8'd67};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd157, 8'd112, 8'd57};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd129, 8'd80, 8'd37};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd135, 8'd90, 8'd57};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd97, 8'd66, 8'd38};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd82, 8'd62, 8'd37};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd103, 8'd73, 8'd37};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd110, 8'd60, 8'd23};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd132, 8'd61, 8'd15};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd167, 8'd89, 8'd25};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd199, 8'd128, 8'd40};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd221, 8'd157, 8'd47};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd240, 8'd176, 8'd50};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd54};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd240, 8'd210, 8'd78};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd242, 8'd211, 8'd84};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd248, 8'd213, 8'd95};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd250, 8'd213, 8'd99};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd253, 8'd209, 8'd100};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd254, 8'd202, 8'd93};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd85};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd77};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd237, 8'd149, 8'd51};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd227, 8'd150, 8'd62};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd206, 8'd134, 8'd60};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd194, 8'd117, 8'd49};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd167, 8'd78, 8'd12};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd153, 8'd59, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd163, 8'd73, 8'd21};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd139, 8'd58, 8'd13};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd121, 8'd99, 8'd101};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd214, 8'd214, 8'd216};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd186, 8'd213, 8'd220};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd148, 8'd187, 8'd202};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd118, 8'd155, 8'd174};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd152, 8'd185, 8'd204};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd142, 8'd176, 8'd188};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd123, 8'd162, 8'd169};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd90, 8'd134, 8'd161};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd97, 8'd137, 8'd162};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd131, 8'd164, 8'd183};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd187, 8'd198, 8'd200};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd175, 8'd174, 8'd170};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd155, 8'd141, 8'd132};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd119, 8'd95, 8'd83};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd127, 8'd62, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd122, 8'd53, 8'd22};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd192, 8'd116, 8'd90};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd155, 8'd80, 8'd57};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd124, 8'd61, 8'd43};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd111, 8'd68, 8'd52};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd142, 8'd120, 8'd106};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd162, 8'd154, 8'd141};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd195, 8'd205, 8'd215};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd179, 8'd199, 8'd206};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd151, 8'd180, 8'd184};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd126, 8'd154, 8'd158};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd122, 8'd139, 8'd147};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd129, 8'd143, 8'd152};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd149, 8'd155};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd115, 8'd149, 8'd151};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd133, 8'd144, 8'd164};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd119, 8'd143, 8'd167};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd90, 8'd130, 8'd155};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd87, 8'd130, 8'd147};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd120, 8'd158, 8'd167};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd121, 8'd155, 8'd164};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd131, 8'd173, 8'd189};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd108, 8'd156, 8'd179};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd144, 8'd172, 8'd196};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd188, 8'd207, 8'd221};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd193, 8'd192, 8'd188};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd136, 8'd98, 8'd79};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd132, 8'd55, 8'd25};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd148, 8'd51, 8'd9};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd161, 8'd64, 8'd11};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd160, 8'd72, 8'd9};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd189, 8'd110, 8'd33};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd201, 8'd125, 8'd41};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd218, 8'd147, 8'd55};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd231, 8'd168, 8'd65};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd238, 8'd182, 8'd73};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd244, 8'd192, 8'd80};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd248, 8'd203, 8'd88};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd252, 8'd209, 8'd94};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd239, 8'd205, 8'd95};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd254, 8'd213, 8'd99};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd95};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd80};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd251, 8'd182, 8'd63};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd238, 8'd165, 8'd54};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd219, 8'd146, 8'd43};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd202, 8'd128, 8'd29};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd152, 8'd85, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd133, 8'd63, 8'd14};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd126, 8'd59, 8'd17};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd122, 8'd66, 8'd31};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd109, 8'd65, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd112, 8'd66, 8'd33};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd138, 8'd74, 8'd46};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd157, 8'd77, 8'd52};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd186, 8'd108, 8'd70};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd198, 8'd138, 8'd76};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd216, 8'd176, 8'd89};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd234, 8'd199, 8'd105};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd249, 8'd204, 8'd119};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd126};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd124};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd254, 8'd213, 8'd121};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd240, 8'd182, 8'd98};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd235, 8'd180, 8'd87};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd224, 8'd171, 8'd67};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd213, 8'd155, 8'd45};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd215, 8'd143, 8'd35};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd222, 8'd127, 8'd33};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd218, 8'd101, 8'd24};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd208, 8'd76, 8'd11};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd190, 8'd19, 8'd2};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd179, 8'd28, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd165, 8'd47, 8'd1};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd148, 8'd60, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd142, 8'd72, 8'd3};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd132, 8'd64, 8'd1};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd129, 8'd53, 8'd1};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd166, 8'd84, 8'd37};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd183, 8'd81, 8'd43};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd197, 8'd103, 8'd51};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd193, 8'd111, 8'd37};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd189, 8'd121, 8'd24};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd204, 8'd146, 8'd36};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd208, 8'd159, 8'd41};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd205, 8'd160, 8'd43};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd214, 8'd169, 8'd54};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd236, 8'd180, 8'd67};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd241, 8'd185, 8'd72};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd248, 8'd195, 8'd83};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd93};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd99};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd100};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd254, 8'd210, 8'd101};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd252, 8'd208, 8'd99};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd237, 8'd231, 8'd109};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd237, 8'd227, 8'd114};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd237, 8'd223, 8'd126};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd240, 8'd219, 8'd136};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd245, 8'd219, 8'd142};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd251, 8'd222, 8'd144};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd144};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd143};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd152};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd168};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd172};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd240, 8'd211, 8'd145};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd215, 8'd163, 8'd90};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd217, 8'd129, 8'd40};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd247, 8'd120, 8'd17};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd126, 8'd13};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd126, 8'd48};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd33};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd231, 8'd165, 8'd9};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd216, 8'd185, 8'd45};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd243, 8'd236, 8'd156};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd72: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd247, 8'd233, 8'd204};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd232, 8'd200, 8'd101};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd235, 8'd170, 8'd6};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd0};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd133, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd111, 8'd41};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd238, 8'd110, 8'd21};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd235, 8'd126, 8'd0};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd234, 8'd107, 8'd36};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd248, 8'd149, 8'd84};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd146};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd181};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd242, 8'd242, 8'd178};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd239, 8'd234, 8'd152};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd249, 8'd227, 8'd126};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd112};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd251, 8'd220, 8'd129};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd251, 8'd220, 8'd127};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd122};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd113};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd104};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd252, 8'd215, 8'd101};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd103};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd108};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd243, 8'd199, 8'd90};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd243, 8'd196, 8'd88};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd240, 8'd192, 8'd84};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd236, 8'd185, 8'd78};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd229, 8'd175, 8'd69};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd221, 8'd162, 8'd58};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd213, 8'd151, 8'd48};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd207, 8'd145, 8'd42};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd212, 8'd125, 8'd28};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd203, 8'd116, 8'd21};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd188, 8'd100, 8'd10};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd168, 8'd81, 8'd1};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd151, 8'd64, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd138, 8'd48, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd127, 8'd38, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd123, 8'd33, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd161, 8'd51, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd170, 8'd55, 8'd11};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd170, 8'd46, 8'd10};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd187, 8'd59, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd208, 8'd88, 8'd35};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd229, 8'd125, 8'd36};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd234, 8'd150, 8'd25};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd248, 8'd179, 8'd26};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd33};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd35};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd252, 8'd154, 8'd43};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd247, 8'd156, 8'd49};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd241, 8'd155, 8'd52};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd236, 8'd154, 8'd52};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd152, 8'd52};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd232, 8'd150, 8'd51};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd235, 8'd151, 8'd52};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd223, 8'd136, 8'd43};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd204, 8'd113, 8'd32};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd186, 8'd93, 8'd26};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd169, 8'd77, 8'd26};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd153, 8'd63, 8'd26};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd138, 8'd53, 8'd24};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd127, 8'd45, 8'd21};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd108, 8'd50, 8'd10};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd115, 8'd63, 8'd16};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd120, 8'd69, 8'd16};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd137, 8'd71, 8'd11};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd182, 8'd95, 8'd26};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd234, 8'd135, 8'd50};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd251, 8'd158, 8'd54};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd40};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd235, 8'd196, 8'd65};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd247, 8'd209, 8'd84};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd252, 8'd217, 8'd101};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd249, 8'd212, 8'd106};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd247, 8'd209, 8'd108};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd253, 8'd211, 8'd111};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd109};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd254, 8'd205, 8'd103};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd249, 8'd200, 8'd98};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd235, 8'd181, 8'd83};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd215, 8'd151, 8'd61};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd184, 8'd113, 8'd31};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd167, 8'd90, 8'd20};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd151, 8'd70, 8'd14};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd162, 8'd81, 8'd34};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd140, 8'd58, 8'd20};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd137, 8'd74, 8'd31};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd217, 8'd185, 8'd162};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd204, 8'd214, 8'd215};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd172, 8'd209, 8'd225};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd146, 8'd187, 8'd205};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd154, 8'd187, 8'd202};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd164, 8'd187, 8'd201};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd168, 8'd190, 8'd204};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd171, 8'd198, 8'd191};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd184, 8'd209, 8'd205};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd203, 8'd223, 8'd224};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd141, 8'd156, 8'd159};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd141, 8'd160, 8'd158};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd187, 8'd206, 8'd200};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd204, 8'd206, 8'd218};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd188, 8'd178, 8'd186};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd181, 8'd153, 8'd152};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd159, 8'd106, 8'd90};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd129, 8'd52, 8'd22};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd117, 8'd25, 8'd0};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd13};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd142, 8'd58, 8'd12};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd191, 8'd118, 8'd73};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd152, 8'd79, 8'd38};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd144, 8'd64, 8'd31};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd136, 8'd57, 8'd27};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd125, 8'd58, 8'd29};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd126, 8'd69, 8'd39};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd144, 8'd126, 8'd114};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd178, 8'd167, 8'd161};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd199, 8'd200, 8'd202};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd181, 8'd191, 8'd200};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd146, 8'd163, 8'd173};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd131, 8'd145, 8'd156};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd134, 8'd143, 8'd152};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd140, 8'd143, 8'd150};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd109, 8'd136, 8'd147};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd104, 8'd133, 8'd141};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd100, 8'd133, 8'd138};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd115, 8'd150, 8'd154};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd147, 8'd185, 8'd188};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd168, 8'd207, 8'd212};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd157, 8'd196, 8'd203};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd132, 8'd169, 8'd178};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd147, 8'd205, 8'd225};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd202, 8'd230, 8'd234};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd215, 8'd190, 8'd170};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd129, 8'd58, 8'd16};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd151, 8'd56, 8'd0};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd144, 8'd49, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd138, 8'd58, 8'd5};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd162, 8'd96, 8'd46};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd188, 8'd107, 8'd44};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd203, 8'd128, 8'd60};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd224, 8'd158, 8'd80};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd238, 8'd182, 8'd95};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd241, 8'd195, 8'd97};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd243, 8'd205, 8'd96};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd247, 8'd212, 8'd96};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd250, 8'd218, 8'd99};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd240, 8'd197, 8'd92};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd251, 8'd214, 8'd97};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd254, 8'd215, 8'd84};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd245, 8'd191, 8'd59};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd237, 8'd161, 8'd41};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd230, 8'd137, 8'd41};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd206, 8'd114, 8'd37};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd181, 8'd96, 8'd32};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd114, 8'd56, 8'd0};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd116, 8'd64, 8'd7};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd124, 8'd75, 8'd34};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd126, 8'd75, 8'd44};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd117, 8'd58, 8'd28};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd117, 8'd43, 8'd4};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd145, 8'd55, 8'd3};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd179, 8'd79, 8'd17};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd179, 8'd89, 8'd26};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd196, 8'd108, 8'd37};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd211, 8'd126, 8'd45};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd222, 8'd139, 8'd47};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd230, 8'd151, 8'd46};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd236, 8'd161, 8'd44};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd234, 8'd160, 8'd37};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd225, 8'd152, 8'd24};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd239, 8'd155, 8'd31};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd245, 8'd157, 8'd24};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd239, 8'd142, 8'd11};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd253, 8'd143, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd249, 8'd122, 8'd45};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd246, 8'd105, 8'd59};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd207, 8'd60, 8'd27};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd166, 8'd15, 8'd0};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd181, 8'd8, 8'd27};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd195, 8'd50, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd195, 8'd74, 8'd21};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd145, 8'd41, 8'd14};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd149, 8'd66, 8'd16};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd122, 8'd41, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd123, 8'd38, 8'd0};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd158, 8'd70, 8'd22};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd164, 8'd88, 8'd26};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd175, 8'd101, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd189, 8'd117, 8'd33};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd201, 8'd133, 8'd36};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd210, 8'd142, 8'd41};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd217, 8'd151, 8'd54};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd226, 8'd159, 8'd68};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd233, 8'd165, 8'd80};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd234, 8'd191, 8'd79};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd234, 8'd192, 8'd80};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd235, 8'd198, 8'd84};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd237, 8'd204, 8'd91};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd243, 8'd210, 8'd97};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd106};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd112};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd115};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd123};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd131};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd140};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd250, 8'd232, 8'd146};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd243, 8'd230, 8'd151};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd243, 8'd229, 8'd156};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd249, 8'd232, 8'd162};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd167};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd163};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd254, 8'd193, 8'd126};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd247, 8'd146, 8'd64};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd242, 8'd108, 8'd11};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd250, 8'd105, 8'd0};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd125, 8'd14};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd248, 8'd143, 8'd28};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd231, 8'd145, 8'd32};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd254, 8'd155, 8'd0};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd235, 8'd155, 8'd18};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd232, 8'd183, 8'd91};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd253, 8'd233, 8'd183};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd73: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd253, 8'd242, 8'd222};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd253, 8'd225, 8'd162};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd245, 8'd190, 8'd74};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd241, 8'd154, 8'd12};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd252, 8'd140, 8'd2};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd141, 8'd20};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd133, 8'd27};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd237, 8'd120, 8'd15};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd246, 8'd113, 8'd12};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd234, 8'd114, 8'd17};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd226, 8'd129, 8'd35};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd230, 8'd160, 8'd74};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd246, 8'd199, 8'd119};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd156};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd170};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd173};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd153};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd252, 8'd230, 8'd144};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd245, 8'd221, 8'd131};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd246, 8'd220, 8'd125};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd124};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd122};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd113};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd252, 8'd214, 8'd107};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd252, 8'd209, 8'd97};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd248, 8'd202, 8'd91};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd241, 8'd190, 8'd81};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd234, 8'd177, 8'd72};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd227, 8'd164, 8'd61};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd221, 8'd153, 8'd52};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd219, 8'd145, 8'd46};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd217, 8'd141, 8'd45};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd212, 8'd122, 8'd36};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd203, 8'd114, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd188, 8'd99, 8'd19};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd169, 8'd81, 8'd10};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd152, 8'd63, 8'd5};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd139, 8'd48, 8'd4};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd128, 8'd37, 8'd6};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd124, 8'd32, 8'd9};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd150, 8'd46, 8'd7};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd171, 8'd57, 8'd23};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd170, 8'd42, 8'd13};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd169, 8'd31, 8'd5};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd188, 8'd54, 8'd17};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd219, 8'd101, 8'd37};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd232, 8'd134, 8'd37};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd239, 8'd156, 8'd34};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd251, 8'd152, 8'd22};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd249, 8'd154, 8'd24};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd247, 8'd158, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd246, 8'd161, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd244, 8'd161, 8'd39};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd243, 8'd160, 8'd40};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd40};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd242, 8'd155, 8'd39};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd228, 8'd135, 8'd32};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd217, 8'd120, 8'd25};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd198, 8'd98, 8'd13};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd180, 8'd77, 8'd8};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd164, 8'd60, 8'd7};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd145, 8'd46, 8'd5};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd128, 8'd33, 8'd1};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd116, 8'd25, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd130, 8'd72, 8'd35};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd121, 8'd72, 8'd31};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd111, 8'd63, 8'd15};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd120, 8'd59, 8'd4};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd162, 8'd81, 8'd16};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd216, 8'd121, 8'd39};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd242, 8'd148, 8'd48};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd239, 8'd154, 8'd38};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd228, 8'd158, 8'd37};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd248, 8'd181, 8'd66};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd98};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd116};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd124};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd123};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd114};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd238, 8'd200, 8'd103};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd237, 8'd191, 8'd103};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd228, 8'd178, 8'd91};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd215, 8'd156, 8'd76};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd194, 8'd128, 8'd54};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd179, 8'd108, 8'd46};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd165, 8'd89, 8'd39};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd175, 8'd97, 8'd58};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd149, 8'd73, 8'd39};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd114, 8'd46, 8'd1};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd184, 8'd147, 8'd121};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd216, 8'd218, 8'd217};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd192, 8'd221, 8'd235};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd158, 8'd194, 8'd210};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd184, 8'd212, 8'd226};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd201, 8'd223, 8'd237};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd178, 8'd197, 8'd212};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd196, 8'd211, 8'd208};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd212, 8'd226, 8'd227};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd226, 8'd237, 8'd241};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd134, 8'd141, 8'd149};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd129, 8'd136, 8'd142};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd182, 8'd192, 8'd193};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd204, 8'd205, 8'd210};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd201, 8'd199, 8'd204};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd179, 8'd167, 8'd169};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd150, 8'd125, 8'd121};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd135, 8'd91, 8'd78};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd126, 8'd61, 8'd39};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd127, 8'd47, 8'd14};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd142, 8'd52, 8'd15};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd154, 8'd56, 8'd17};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd142, 8'd58, 8'd14};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd191, 8'd116, 8'd74};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd155, 8'd77, 8'd38};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd147, 8'd63, 8'd29};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd143, 8'd56, 8'd26};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd132, 8'd56, 8'd24};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd132, 8'd68, 8'd33};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd113, 8'd78, 8'd59};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd143, 8'd117, 8'd104};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd172, 8'd161, 8'd157};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd180, 8'd181, 8'd185};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd169, 8'd179, 8'd188};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd157, 8'd170, 8'd179};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd153, 8'd163, 8'd172};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd151, 8'd160, 8'd167};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd109, 8'd126, 8'd142};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd102, 8'd121, 8'd135};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd99, 8'd123, 8'd135};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd111, 8'd138, 8'd147};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd130, 8'd159, 8'd167};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd147, 8'd174, 8'd183};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd156, 8'd183, 8'd194};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd161, 8'd185, 8'd197};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd186, 8'd224, 8'd235};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd226, 8'd235, 8'd234};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd185, 8'd150, 8'd130};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd132, 8'd57, 8'd18};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd7};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd12};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd137, 8'd59, 8'd20};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd143, 8'd79, 8'd44};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd180, 8'd105, 8'd50};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd194, 8'd124, 8'd64};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd215, 8'd150, 8'd84};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd230, 8'd173, 8'd96};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd237, 8'd187, 8'd100};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd241, 8'd197, 8'd102};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd247, 8'd205, 8'd103};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd106};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd107};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd88};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd239, 8'd184, 8'd58};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd228, 8'd160, 8'd33};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd236, 8'd146, 8'd34};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd236, 8'd135, 8'd45};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd212, 8'd113, 8'd45};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd180, 8'd89, 8'd32};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd117, 8'd61, 8'd4};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd121, 8'd67, 8'd20};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd126, 8'd73, 8'd39};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd123, 8'd67, 8'd40};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd116, 8'd52, 8'd24};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd124, 8'd46, 8'd7};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd151, 8'd60, 8'd5};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd179, 8'd80, 8'd13};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd194, 8'd94, 8'd16};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd210, 8'd111, 8'd26};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd224, 8'd130, 8'd34};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd234, 8'd143, 8'd36};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd243, 8'd154, 8'd36};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd248, 8'd163, 8'd36};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd245, 8'd161, 8'd29};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd236, 8'd154, 8'd19};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd244, 8'd161, 8'd31};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd250, 8'd161, 8'd31};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd242, 8'd142, 8'd20};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd245, 8'd128, 8'd33};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd224, 8'd92, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd216, 8'd72, 8'd35};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd190, 8'd39, 8'd8};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd170, 8'd17, 8'd0};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd179, 8'd22, 8'd13};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd228, 8'd96, 8'd24};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd232, 8'd118, 8'd58};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd141, 8'd41, 8'd18};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd127, 8'd42, 8'd1};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd119, 8'd38, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd133, 8'd46, 8'd3};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd157, 8'd67, 8'd14};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd171, 8'd81, 8'd19};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd180, 8'd93, 8'd22};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd193, 8'd108, 8'd25};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd202, 8'd122, 8'd27};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd206, 8'd131, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd213, 8'd139, 8'd40};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd221, 8'd146, 8'd53};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd227, 8'd153, 8'd66};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd221, 8'd163, 8'd55};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd226, 8'd174, 8'd64};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd236, 8'd193, 8'd81};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd244, 8'd211, 8'd98};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd251, 8'd224, 8'd111};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd253, 8'd230, 8'd118};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd252, 8'd230, 8'd119};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd251, 8'd229, 8'd118};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd121};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd243, 8'd224, 8'd122};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd245, 8'd225, 8'd130};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd254, 8'd230, 8'd142};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd151};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd152};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd140};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd130};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd226, 8'd142, 8'd78};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd221, 8'd127, 8'd57};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd232, 8'd121, 8'd39};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd251, 8'd127, 8'd31};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd128, 8'd15};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd249, 8'd127, 8'd0};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd6};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd27};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd239, 8'd157, 8'd29};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd244, 8'd179, 8'd75};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd253, 8'd214, 8'd147};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd217};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd74: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd168};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd237, 8'd181, 8'd72};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd236, 8'd162, 8'd5};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd0};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd19};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd252, 8'd129, 8'd35};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd241, 8'd126, 8'd7};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd250, 8'd130, 8'd8};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd253, 8'd127, 8'd7};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd242, 8'd118, 8'd4};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd223, 8'd115, 8'd14};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd217, 8'd136, 8'd54};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd229, 8'd175, 8'd111};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd243, 8'd208, 8'd154};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd153};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd150};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd145};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd254, 8'd224, 8'd138};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd129};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd251, 8'd218, 8'd125};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd253, 8'd219, 8'd122};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd254, 8'd220, 8'd123};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd252, 8'd215, 8'd100};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd249, 8'd208, 8'd94};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd244, 8'd194, 8'd83};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd235, 8'd177, 8'd70};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd227, 8'd158, 8'd57};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd220, 8'd142, 8'd44};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd214, 8'd129, 8'd36};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd212, 8'd123, 8'd31};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd211, 8'd120, 8'd41};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd203, 8'd111, 8'd34};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd189, 8'd98, 8'd25};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd173, 8'd81, 8'd18};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd155, 8'd63, 8'd12};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd140, 8'd48, 8'd11};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd131, 8'd37, 8'd12};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd126, 8'd30, 8'd14};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd127, 8'd31, 8'd6};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd176, 8'd67, 8'd38};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd192, 8'd61, 8'd31};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd169, 8'd20, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd169, 8'd17, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd196, 8'd56, 8'd23};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd220, 8'd99, 8'd42};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd232, 8'd127, 8'd46};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd237, 8'd150, 8'd11};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd237, 8'd154, 8'd14};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd241, 8'd160, 8'd19};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd244, 8'd164, 8'd23};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd248, 8'd167, 8'd26};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd249, 8'd166, 8'd26};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd253, 8'd163, 8'd27};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd253, 8'd161, 8'd26};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd252, 8'd150, 8'd40};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd242, 8'd136, 8'd34};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd224, 8'd114, 8'd25};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd207, 8'd95, 8'd21};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd190, 8'd77, 8'd17};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd169, 8'd61, 8'd14};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd149, 8'd45, 8'd8};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd136, 8'd36, 8'd4};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd113, 8'd53, 8'd25};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd114, 8'd65, 8'd33};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd112, 8'd68, 8'd29};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd113, 8'd59, 8'd13};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd133, 8'd61, 8'd3};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd176, 8'd88, 8'd14};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd218, 8'd127, 8'd34};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd241, 8'd156, 8'd47};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd38};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd54};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd69};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd243, 8'd175, 8'd76};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd237, 8'd183, 8'd87};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd244, 8'd200, 8'd105};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd118};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd254, 8'd218, 8'd124};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd243, 8'd197, 8'd122};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd235, 8'd185, 8'd112};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd218, 8'd161, 8'd92};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd187, 8'd121, 8'd60};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd162, 8'd91, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd144, 8'd71, 8'd28};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd164, 8'd90, 8'd55};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd150, 8'd76, 8'd47};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd150, 8'd77, 8'd32};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd147, 8'd103, 8'd76};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd210, 8'd205, 8'd202};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd232, 8'd250, 8'd255};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd197, 8'd220, 8'd234};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd205, 8'd219};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd214, 8'd230, 8'd245};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd221, 8'd237, 8'd253};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd233, 8'd238, 8'd241};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd242, 8'd247, 8'd251};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd255};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd235, 8'd237, 8'd249};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd200, 8'd200, 8'd212};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd188, 8'd186, 8'd197};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd205, 8'd202, 8'd209};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd219, 8'd217, 8'd222};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd178, 8'd166, 8'd168};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd162, 8'd141, 8'd136};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd129, 8'd93, 8'd81};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd110, 8'd58, 8'd36};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd121, 8'd52, 8'd23};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd130, 8'd50, 8'd17};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd134, 8'd48, 8'd13};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd146, 8'd56, 8'd21};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd154, 8'd57, 8'd24};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd142, 8'd57, 8'd20};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd192, 8'd114, 8'd75};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd157, 8'd75, 8'd37};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd154, 8'd61, 8'd27};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd22};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd142, 8'd54, 8'd18};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd142, 8'd63, 8'd24};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd115, 8'd54, 8'd25};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd110, 8'd58, 8'd36};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd117, 8'd83, 8'd71};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd144, 8'd129, 8'd126};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd174, 8'd173, 8'd178};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd185, 8'd192, 8'd200};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd175, 8'd188, 8'd196};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd164, 8'd177, 8'd183};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd113, 8'd121, 8'd140};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd104, 8'd115, 8'd133};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd104, 8'd121, 8'd137};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd119, 8'd138, 8'd153};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd129, 8'd148, 8'd162};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd134, 8'd152, 8'd164};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd148, 8'd162, 8'd175};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd166, 8'd176, 8'd188};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd207, 8'd225, 8'd227};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd237, 8'd230, 8'd222};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd163, 8'd121, 8'd99};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd148, 8'd74, 8'd39};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd156, 8'd63, 8'd22};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd166, 8'd72, 8'd34};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd150, 8'd67, 8'd33};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd151, 8'd77, 8'd48};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd173, 8'd101, 8'd53};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd185, 8'd115, 8'd64};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd202, 8'd133, 8'd76};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd215, 8'd150, 8'd86};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd225, 8'd161, 8'd90};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd230, 8'd168, 8'd91};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd234, 8'd176, 8'd92};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd238, 8'd182, 8'd95};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd235, 8'd153, 8'd51};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd230, 8'd157, 8'd46};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd228, 8'd158, 8'd37};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd234, 8'd153, 8'd35};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd242, 8'd145, 8'd42};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd225, 8'd120, 8'd39};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd175, 8'd75, 8'd13};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd126, 8'd36, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd123, 8'd66, 8'd23};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd128, 8'd72, 8'd37};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd128, 8'd71, 8'd44};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd118, 8'd56, 8'd33};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd116, 8'd45, 8'd15};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd134, 8'd52, 8'd5};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd163, 8'd69, 8'd7};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd184, 8'd84, 8'd9};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd210, 8'd103, 8'd5};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd226, 8'd121, 8'd16};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd239, 8'd138, 8'd24};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd248, 8'd148, 8'd24};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd28};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd24};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd247, 8'd153, 8'd17};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd239, 8'd157, 8'd22};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd245, 8'd153, 8'd28};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd236, 8'd129, 8'd25};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd224, 8'd99, 8'd32};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd196, 8'd54, 8'd18};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd187, 8'd37, 8'd13};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd180, 8'd27, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd191, 8'd38, 8'd0};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd223, 8'd93, 8'd43};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd47};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd227, 8'd126, 8'd56};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd112, 8'd17, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd110, 8'd25, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd129, 8'd45, 8'd1};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd148, 8'd57, 8'd13};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd154, 8'd62, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd183, 8'd81, 8'd17};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd192, 8'd91, 8'd19};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd202, 8'd107, 8'd23};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd208, 8'd119, 8'd25};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd211, 8'd127, 8'd28};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd215, 8'd135, 8'd36};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd221, 8'd142, 8'd47};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd225, 8'd149, 8'd55};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd235, 8'd167, 8'd58};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd238, 8'd178, 8'd68};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd240, 8'd192, 8'd81};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd243, 8'd207, 8'd95};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd243, 8'd220, 8'd108};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd241, 8'd225, 8'd114};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd239, 8'd227, 8'd117};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd237, 8'd226, 8'd118};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd234, 8'd219, 8'd116};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd247, 8'd227, 8'd128};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd140};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd139};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd117};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd242, 8'd160, 8'd78};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd219, 8'd120, 8'd37};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd204, 8'd95, 8'd13};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd229, 8'd96, 8'd17};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd237, 8'd108, 8'd24};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd244, 8'd121, 8'd27};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd248, 8'd133, 8'd24};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd251, 8'd143, 8'd17};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd254, 8'd152, 8'd8};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd0};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd0};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd231, 8'd180, 8'd99};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd154};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd215};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd75: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd253, 8'd227, 8'd166};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd241, 8'd199, 8'd78};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd237, 8'd172, 8'd16};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd248, 8'd157, 8'd8};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd26};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd238, 8'd154, 8'd29};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd244, 8'd145, 8'd18};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd251, 8'd129, 8'd4};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd252, 8'd113, 8'd0};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd250, 8'd106, 8'd0};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd244, 8'd111, 8'd10};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd241, 8'd123, 8'd33};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd241, 8'd135, 8'd51};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd224, 8'd155, 8'd78};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd241, 8'd174, 8'd96};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd120};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd134};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd134};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd126};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd252, 8'd218, 8'd120};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd115};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd240, 8'd208, 8'd87};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd238, 8'd202, 8'd82};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd234, 8'd189, 8'd74};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd229, 8'd173, 8'd64};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd226, 8'd159, 8'd55};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd224, 8'd146, 8'd48};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd225, 8'd138, 8'd45};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd224, 8'd133, 8'd42};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd209, 8'd117, 8'd32};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd202, 8'd111, 8'd28};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd190, 8'd98, 8'd21};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd175, 8'd84, 8'd14};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd160, 8'd67, 8'd10};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd144, 8'd51, 8'd8};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd133, 8'd39, 8'd11};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd127, 8'd32, 8'd10};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd104, 8'd16, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd183, 8'd81, 8'd43};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd232, 8'd108, 8'd57};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd201, 8'd54, 8'd11};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd175, 8'd15, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd171, 8'd14, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd199, 8'd59, 8'd26};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd226, 8'd96, 8'd47};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd219, 8'd135, 8'd13};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd141, 8'd15};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd232, 8'd151, 8'd18};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd240, 8'd160, 8'd21};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd248, 8'd165, 8'd23};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd25};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd23};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd25};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd38};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd247, 8'd146, 8'd32};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd233, 8'd127, 8'd25};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd217, 8'd109, 8'd21};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd199, 8'd91, 8'd19};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd177, 8'd72, 8'd14};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd154, 8'd54, 8'd4};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd139, 8'd42, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd94, 8'd28, 8'd6};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd106, 8'd52, 8'd26};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd116, 8'd75, 8'd45};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd119, 8'd74, 8'd35};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd121, 8'd57, 8'd9};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd142, 8'd61, 8'd0};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd182, 8'd96, 8'd11};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd217, 8'd133, 8'd34};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd246, 8'd140, 8'd20};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd252, 8'd153, 8'd34};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd48};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd239, 8'd163, 8'd53};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd233, 8'd166, 8'd62};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd238, 8'd176, 8'd77};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd241, 8'd182, 8'd88};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd239, 8'd183, 8'd90};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd235, 8'd178, 8'd109};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd227, 8'd166, 8'd99};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd216, 8'd148, 8'd85};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd192, 8'd120, 8'd61};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd179, 8'd103, 8'd51};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd165, 8'd88, 8'd46};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd178, 8'd102, 8'd68};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd156, 8'd81, 8'd50};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd121, 8'd53, 8'd8};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd136, 8'd92, 8'd67};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd222, 8'd211, 8'd207};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd232, 8'd240, 8'd251};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd213, 8'd225, 8'd237};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd219, 8'd229, 8'd239};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd236, 8'd248, 8'd255};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd223, 8'd237, 8'd250};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd228, 8'd233, 8'd236};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd230, 8'd235, 8'd239};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd238, 8'd242, 8'd251};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd245, 8'd248, 8'd255};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd240, 8'd240, 8'd250};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd223, 8'd218, 8'd225};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd195, 8'd186, 8'd191};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd171, 8'd159, 8'd161};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd154, 8'd125, 8'd119};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd130, 8'd88, 8'd74};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd100, 8'd40, 8'd14};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd105, 8'd27, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd145, 8'd53, 8'd12};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd163, 8'd67, 8'd25};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd150, 8'd56, 8'd18};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd138, 8'd48, 8'd13};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd157, 8'd59, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd144, 8'd55, 8'd21};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd193, 8'd111, 8'd73};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd161, 8'd73, 8'd35};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd161, 8'd61, 8'd25};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd162, 8'd55, 8'd19};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd150, 8'd51, 8'd10};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd150, 8'd59, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd146, 8'd61, 8'd22};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd110, 8'd35, 8'd3};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd86, 8'd28, 8'd8};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd103, 8'd65, 8'd56};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd140, 8'd120, 8'd121};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd165, 8'd160, 8'd164};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd175, 8'd180, 8'd183};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd179, 8'd189, 8'd190};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd141, 8'd148, 8'd164};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd128, 8'd140, 8'd156};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd120, 8'd137, 8'd153};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd122, 8'd145, 8'd159};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd129, 8'd152, 8'd166};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd133, 8'd153, 8'd164};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd138, 8'd152, 8'd163};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd146, 8'd154, 8'd165};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd171, 8'd187, 8'd186};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd196, 8'd193, 8'd184};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd153, 8'd121, 8'd98};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd158, 8'd95, 8'd60};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd159, 8'd76, 8'd32};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd171, 8'd79, 8'd32};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd158, 8'd66, 8'd19};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd169, 8'd81, 8'd35};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd167, 8'd91, 8'd42};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd174, 8'd96, 8'd47};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd185, 8'd104, 8'd51};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd196, 8'd111, 8'd54};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd204, 8'd119, 8'd55};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd209, 8'd125, 8'd55};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd212, 8'd130, 8'd56};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd215, 8'd133, 8'd57};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd220, 8'd131, 8'd31};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd225, 8'd144, 8'd37};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd230, 8'd155, 8'd40};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd230, 8'd150, 8'd39};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd221, 8'd128, 8'd33};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd195, 8'd99, 8'd23};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd156, 8'd70, 8'd13};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd125, 8'd51, 8'd2};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd127, 8'd72, 8'd42};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd133, 8'd76, 8'd49};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd128, 8'd66, 8'd45};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd116, 8'd45, 8'd23};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd121, 8'd41, 8'd8};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd146, 8'd59, 8'd6};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd174, 8'd80, 8'd8};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd189, 8'd90, 8'd5};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd220, 8'd115, 8'd8};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd234, 8'd130, 8'd17};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd246, 8'd146, 8'd22};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd252, 8'd155, 8'd24};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd26};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd33};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd244, 8'd151, 8'd22};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd227, 8'd140, 8'd11};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd225, 8'd128, 8'd15};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd215, 8'd98, 8'd18};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd204, 8'd66, 8'd27};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd180, 8'd28, 8'd17};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd179, 8'd22, 8'd13};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd184, 8'd31, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd224, 8'd75, 8'd19};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd69};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd39};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd201, 8'd112, 8'd32};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd96, 8'd7, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd116, 8'd29, 8'd10};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd137, 8'd49, 8'd13};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd147, 8'd54, 8'd11};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd152, 8'd58, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd181, 8'd78, 8'd9};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd190, 8'd90, 8'd14};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd201, 8'd105, 8'd19};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd207, 8'd119, 8'd22};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd210, 8'd127, 8'd25};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd214, 8'd135, 8'd32};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd219, 8'd144, 8'd42};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd224, 8'd151, 8'd49};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd234, 8'd173, 8'd58};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd238, 8'd181, 8'd66};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd243, 8'd196, 8'd82};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd210, 8'd97};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd254, 8'd220, 8'd112};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd120};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd123};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd125};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd135};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd120};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd245, 8'd178, 8'd91};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd226, 8'd142, 8'd56};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd216, 8'd115, 8'd27};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd225, 8'd108, 8'd15};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd247, 8'd117, 8'd21};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd128, 8'd29};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd118, 8'd13};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd135, 8'd21};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd143, 8'd16};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd249, 8'd144, 8'd3};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd243, 8'd151, 8'd6};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd247, 8'd166, 8'd23};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd33};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd228, 8'd161, 8'd31};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd240, 8'd219, 8'd176};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd215};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd76: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd187};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd242, 8'd195, 8'd103};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd239, 8'd170, 8'd33};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd249, 8'd166, 8'd2};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd254, 8'd163, 8'd20};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd249, 8'd151, 8'd14};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd249, 8'd140, 8'd13};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd138, 8'd21};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd141, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd136, 8'd28};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd121, 8'd15};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd107, 8'd0};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd234, 8'd109, 8'd25};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd233, 8'd115, 8'd28};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd235, 8'd130, 8'd39};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd244, 8'd154, 8'd58};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd80};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd95};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd100};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd252, 8'd212, 8'd99};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd97};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd251, 8'd211, 8'd89};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd241, 8'd194, 8'd78};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd232, 8'd176, 8'd65};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd226, 8'd159, 8'd55};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd222, 8'd146, 8'd48};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd221, 8'd138, 8'd44};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd222, 8'd134, 8'd44};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd207, 8'd117, 8'd20};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd202, 8'd112, 8'd16};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd192, 8'd101, 8'd12};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd178, 8'd87, 8'd6};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd163, 8'd72, 8'd2};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd149, 8'd55, 8'd1};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd136, 8'd43, 8'd2};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd130, 8'd36, 8'd2};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd102, 8'd15, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd184, 8'd90, 8'd36};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd65};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd242, 8'd111, 8'd33};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd209, 8'd58, 8'd13};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd166, 8'd7, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd182, 8'd27, 8'd5};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd210, 8'd60, 8'd27};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd203, 8'd107, 8'd21};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd210, 8'd115, 8'd23};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd222, 8'd131, 8'd26};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd233, 8'd147, 8'd28};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd245, 8'd156, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd253, 8'd161, 8'd28};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd246, 8'd158, 8'd25};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd239, 8'd147, 8'd22};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd227, 8'd131, 8'd18};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd213, 8'd115, 8'd16};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd197, 8'd98, 8'd15};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd173, 8'd79, 8'd9};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd148, 8'd58, 8'd0};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd133, 8'd44, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd112, 8'd31, 8'd10};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd108, 8'd46, 8'd23};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd114, 8'd70, 8'd43};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd125, 8'd81, 8'd52};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd130, 8'd72, 8'd34};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd135, 8'd62, 8'd7};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd160, 8'd81, 8'd6};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd190, 8'd110, 8'd21};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd231, 8'd148, 8'd18};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd244, 8'd162, 8'd34};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd249, 8'd171, 8'd45};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd242, 8'd168, 8'd47};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd235, 8'd159, 8'd47};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd233, 8'd154, 8'd51};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd229, 8'd146, 8'd52};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd224, 8'd136, 8'd47};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd202, 8'd129, 8'd61};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd191, 8'd116, 8'd49};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd183, 8'd103, 8'd40};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd173, 8'd93, 8'd34};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd173, 8'd93, 8'd40};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd159, 8'd82, 8'd38};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd158, 8'd84, 8'd49};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd121, 8'd50, 8'd18};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd141, 8'd83, 8'd45};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd156, 8'd120, 8'd98};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd216, 8'd204, 8'd204};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd219, 8'd223, 8'd234};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd232, 8'd239, 8'd249};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd235, 8'd240, 8'd246};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd212, 8'd221, 8'd228};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd179, 8'd192, 8'd201};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd219, 8'd229, 8'd230};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd222, 8'd234, 8'd234};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd223, 8'd234, 8'd236};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd219, 8'd227, 8'd229};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd209, 8'd209, 8'd209};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd183, 8'd173, 8'd171};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd153, 8'd134, 8'd127};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd134, 8'd110, 8'd100};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd128, 8'd77, 8'd60};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd121, 8'd59, 8'd36};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd111, 8'd32, 8'd0};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd124, 8'd31, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd159, 8'd57, 8'd9};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd170, 8'd67, 8'd22};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd156, 8'd58, 8'd19};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd147, 8'd53, 8'd17};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd160, 8'd61, 8'd32};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd145, 8'd55, 8'd21};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd193, 8'd109, 8'd72};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd163, 8'd71, 8'd32};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd168, 8'd62, 8'd23};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd169, 8'd57, 8'd19};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd157, 8'd50, 8'd8};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd152, 8'd56, 8'd8};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd157, 8'd59, 8'd12};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd130, 8'd41, 8'd1};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd105, 8'd29, 8'd3};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd97, 8'd38, 8'd24};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd101, 8'd60, 8'd54};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd116, 8'd91, 8'd86};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd146, 8'd133, 8'd125};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd175, 8'd166, 8'd157};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd173, 8'd178, 8'd182};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd164, 8'd175, 8'd181};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd145, 8'd165, 8'd174};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd125, 8'd153, 8'd164};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd119, 8'd151, 8'd162};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd127, 8'd156, 8'd164};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd135, 8'd155, 8'd162};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd136, 8'd151, 8'd158};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd124, 8'd154, 8'd156};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd137, 8'd154, 8'd148};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd148, 8'd139, 8'd122};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd151, 8'd115, 8'd83};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd162, 8'd101, 8'd54};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd172, 8'd92, 8'd33};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd155, 8'd63, 8'd0};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd170, 8'd73, 8'd2};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd154, 8'd73, 8'd17};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd158, 8'd72, 8'd15};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd165, 8'd70, 8'd14};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd173, 8'd73, 8'd13};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd183, 8'd79, 8'd16};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd191, 8'd88, 8'd21};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd195, 8'd94, 8'd22};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd195, 8'd97, 8'd22};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd197, 8'd113, 8'd17};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd200, 8'd127, 8'd25};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd205, 8'd138, 8'd33};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd200, 8'd131, 8'd28};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd183, 8'd103, 8'd16};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd155, 8'd76, 8'd7};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd133, 8'd66, 8'd11};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd121, 8'd67, 8'd20};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd128, 8'd76, 8'd52};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd131, 8'd73, 8'd51};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd126, 8'd58, 8'd37};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd119, 8'd39, 8'd14};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd131, 8'd41, 8'd4};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd161, 8'd67, 8'd6};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd187, 8'd90, 8'd9};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd198, 8'd99, 8'd6};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd222, 8'd124, 8'd17};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd235, 8'd139, 8'd26};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd246, 8'd152, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd249, 8'd158, 8'd28};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd251, 8'd160, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd250, 8'd160, 8'd37};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd241, 8'd151, 8'd37};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd229, 8'd138, 8'd31};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd219, 8'd121, 8'd14};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd209, 8'd98, 8'd9};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd198, 8'd67, 8'd11};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd191, 8'd41, 8'd26};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd177, 8'd18, 8'd23};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd180, 8'd22, 8'd19};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd186, 8'd38, 8'd2};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd244, 8'd102, 8'd38};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd248, 8'd160, 8'd50};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd243, 8'd163, 8'd22};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd199, 8'd117, 8'd31};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd109, 8'd19, 8'd8};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd124, 8'd35, 8'd21};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd129, 8'd38, 8'd7};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd138, 8'd42, 8'd0};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd154, 8'd57, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd172, 8'd76, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd180, 8'd87, 8'd7};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd193, 8'd103, 8'd15};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd201, 8'd117, 8'd21};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd205, 8'd126, 8'd25};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd212, 8'd135, 8'd31};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd217, 8'd144, 8'd39};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd224, 8'd151, 8'd46};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd238, 8'd183, 8'd66};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd247, 8'd192, 8'd75};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd90};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd101};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd104};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd99};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd89};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd251, 8'd174, 8'd82};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd226, 8'd124, 8'd40};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd222, 8'd116, 8'd32};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd222, 8'd107, 8'd24};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd229, 8'd107, 8'd21};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd243, 8'd114, 8'd20};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd122, 8'd17};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd125, 8'd10};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd124, 8'd4};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd19};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd253, 8'd146, 8'd4};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd0};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd0};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd243, 8'd163, 8'd16};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd224, 8'd169, 8'd52};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd229, 8'd198, 8'd115};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd248, 8'd232, 8'd170};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd77: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd207};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd246, 8'd202, 8'd107};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd230, 8'd179, 8'd28};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd3};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd15};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd28};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd34};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd247, 8'd146, 8'd32};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd245, 8'd135, 8'd24};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd128, 8'd19};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd127, 8'd18};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd117, 8'd19};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd253, 8'd111, 8'd11};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd237, 8'd105, 8'd4};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd225, 8'd108, 8'd2};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd222, 8'd120, 8'd10};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd227, 8'd140, 8'd27};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd236, 8'd159, 8'd43};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd242, 8'd171, 8'd55};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd72};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd189, 8'd74};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd74};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd252, 8'd178, 8'd71};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd244, 8'd165, 8'd64};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd230, 8'd147, 8'd51};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd218, 8'd130, 8'd40};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd209, 8'd121, 8'd32};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd206, 8'd114, 8'd13};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd202, 8'd110, 8'd11};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd193, 8'd103, 8'd7};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd181, 8'd89, 8'd2};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd166, 8'd74, 8'd1};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd151, 8'd58, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd139, 8'd44, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd131, 8'd37, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd115, 8'd22, 8'd7};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd177, 8'd88, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd48};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd36};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd237, 8'd113, 8'd41};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd178, 8'd30, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd177, 8'd16, 8'd0};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd197, 8'd29, 8'd3};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd192, 8'd71, 8'd26};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd199, 8'd84, 8'd27};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd212, 8'd104, 8'd29};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd225, 8'd125, 8'd29};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd237, 8'd141, 8'd29};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd245, 8'd150, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd250, 8'd152, 8'd29};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd251, 8'd151, 8'd29};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd247, 8'd159, 8'd23};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd243, 8'd152, 8'd20};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd234, 8'd141, 8'd22};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd224, 8'd127, 8'd24};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd207, 8'd112, 8'd22};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd185, 8'd92, 8'd15};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd159, 8'd70, 8'd4};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd141, 8'd55, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd125, 8'd25, 8'd1};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd112, 8'd34, 8'd11};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd112, 8'd60, 8'd36};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd126, 8'd84, 8'd59};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd132, 8'd82, 8'd49};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd138, 8'd72, 8'd24};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd167, 8'd93, 8'd28};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd205, 8'd132, 8'd53};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd235, 8'd170, 8'd50};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd241, 8'd177, 8'd54};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd237, 8'd172, 8'd52};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd222, 8'd155, 8'd38};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd214, 8'd141, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd218, 8'd134, 8'd35};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd223, 8'd129, 8'd41};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd223, 8'd122, 8'd40};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd208, 8'd124, 8'd60};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd199, 8'd115, 8'd51};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd181, 8'd99, 8'd39};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd156, 8'd77, 8'd21};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd144, 8'd72, 8'd24};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd143, 8'd78, 8'd40};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd173, 8'd116, 8'd86};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd166, 8'd112, 8'd88};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd195, 8'd158, 8'd131};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd223, 8'd201, 8'd188};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd251, 8'd249, 8'd254};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd229, 8'd235, 8'd247};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd199, 8'd202, 8'd211};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd174, 8'd175, 8'd179};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd189, 8'd197, 8'd199};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd230, 8'd244, 8'd247};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd229, 8'd238, 8'd237};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd229, 8'd240, 8'd236};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd214, 8'd223, 8'd218};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd193, 8'd194, 8'd188};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd149};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd146, 8'd119, 8'd102};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd125, 8'd83, 8'd61};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd122, 8'd70, 8'd46};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd132, 8'd56, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd128, 8'd49, 8'd19};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd120, 8'd31, 8'd0};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd129, 8'd33, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd153, 8'd54, 8'd12};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd164, 8'd63, 8'd21};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd158, 8'd56, 8'd16};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd156, 8'd57, 8'd18};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd163, 8'd63, 8'd29};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd147, 8'd55, 8'd18};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd192, 8'd107, 8'd66};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd162, 8'd70, 8'd29};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd23};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd171, 8'd59, 8'd19};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd157, 8'd52, 8'd7};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd7};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd4};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd140, 8'd47, 8'd4};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd127, 8'd40, 8'd12};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd113, 8'd38, 8'd17};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd104, 8'd41, 8'd26};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd106, 8'd54, 8'd40};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd121, 8'd80, 8'd60};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd139, 8'd103, 8'd79};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd162, 8'd152, 8'd143};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd170, 8'd169, 8'd165};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd164, 8'd178, 8'd179};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd144, 8'd169, 8'd174};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd129, 8'd159, 8'd169};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd131, 8'd160, 8'd168};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd135, 8'd158, 8'd164};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd134, 8'd152, 8'd156};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd127, 8'd160, 8'd169};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd124, 8'd149, 8'd153};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd152, 8'd165, 8'd158};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd147, 8'd140, 8'd122};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd170, 8'd141, 8'd107};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd179, 8'd129, 8'd78};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd162, 8'd94, 8'd31};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd162, 8'd84, 8'd12};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd150, 8'd71, 8'd12};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd149, 8'd65, 8'd5};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd151, 8'd56, 8'd0};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd159, 8'd56, 8'd0};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd1};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd179, 8'd74, 8'd8};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd181, 8'd83, 8'd12};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd183, 8'd87, 8'd13};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd192, 8'd111, 8'd29};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd192, 8'd122, 8'd34};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd198, 8'd137, 8'd44};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd207, 8'd143, 8'd55};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd197, 8'd125, 8'd49};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd167, 8'd97, 8'd35};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd138, 8'd83, 8'd29};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd123, 8'd81, 8'd33};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd127, 8'd80, 8'd52};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd124, 8'd68, 8'd43};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd121, 8'd49, 8'd24};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd125, 8'd38, 8'd8};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd146, 8'd48, 8'd3};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd176, 8'd74, 8'd8};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd198, 8'd98, 8'd12};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd207, 8'd109, 8'd8};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd227, 8'd128, 8'd24};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd238, 8'd142, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd246, 8'd151, 8'd31};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd244, 8'd152, 8'd27};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd241, 8'd151, 8'd29};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd237, 8'd145, 8'd36};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd225, 8'd132, 8'd37};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd212, 8'd118, 8'd31};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd217, 8'd101, 8'd28};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd200, 8'd71, 8'd13};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd190, 8'd46, 8'd12};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd188, 8'd29, 8'd26};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd181, 8'd17, 8'd28};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd179, 8'd21, 8'd18};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd175, 8'd33, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd243, 8'd112, 8'd40};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd238, 8'd154, 8'd42};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd240, 8'd165, 8'd20};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd200, 8'd119, 8'd28};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd105, 8'd13, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd116, 8'd24, 8'd9};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd128, 8'd35, 8'd4};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd142, 8'd44, 8'd7};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd159, 8'd61, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd180, 8'd87, 8'd9};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd189, 8'd96, 8'd16};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd202, 8'd110, 8'd25};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd210, 8'd121, 8'd31};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd215, 8'd128, 8'd33};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd221, 8'd135, 8'd36};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd229, 8'd143, 8'd42};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd233, 8'd150, 8'd46};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd247, 8'd175, 8'd64};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd249, 8'd176, 8'd65};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd251, 8'd175, 8'd65};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd169, 8'd62};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd247, 8'd155, 8'd52};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd240, 8'd138, 8'd40};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd232, 8'd119, 8'd25};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd227, 8'd108, 8'd16};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd117, 8'd26};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd115, 8'd25};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd253, 8'd115, 8'd24};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd121, 8'd22};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd130, 8'd22};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd139, 8'd19};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd17};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd14};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd242, 8'd161, 8'd17};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd242, 8'd158, 8'd8};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd6};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd243, 8'd163, 8'd22};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd239, 8'd179, 8'd65};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd236, 8'd204, 8'd131};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd240, 8'd237, 8'd204};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd78: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd196};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd241, 8'd214, 8'd135};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd74};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd251, 8'd167, 8'd53};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd235, 8'd153, 8'd27};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd231, 8'd149, 8'd13};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd239, 8'd153, 8'd14};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd248, 8'd155, 8'd24};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd150, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd249, 8'd143, 8'd31};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd124, 8'd10};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd131, 8'd17};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd137, 8'd24};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd132, 8'd22};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd245, 8'd120, 8'd12};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd232, 8'd111, 8'd4};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd226, 8'd108, 8'd2};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd227, 8'd108, 8'd4};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd231, 8'd122, 8'd17};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd236, 8'd127, 8'd24};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd243, 8'd135, 8'd34};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd248, 8'd141, 8'd45};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd244, 8'd141, 8'd48};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd236, 8'd135, 8'd45};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd227, 8'd127, 8'd41};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd221, 8'd121, 8'd36};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd205, 8'd112, 8'd17};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd202, 8'd109, 8'd16};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd195, 8'd101, 8'd13};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd183, 8'd90, 8'd12};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd168, 8'd75, 8'd8};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd154, 8'd58, 8'd7};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd141, 8'd45, 8'd5};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd133, 8'd36, 8'd4};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd119, 8'd14, 8'd18};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd167, 8'd79, 8'd15};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd235, 8'd162, 8'd33};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd238, 8'd165, 8'd26};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd238, 8'd140, 8'd51};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd181, 8'd48, 8'd15};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd183, 8'd21, 8'd10};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd199, 8'd19, 8'd5};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd184, 8'd39, 8'd22};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd192, 8'd53, 8'd22};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd204, 8'd79, 8'd21};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd217, 8'd107, 8'd22};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd128, 8'd22};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd235, 8'd140, 8'd22};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd237, 8'd145, 8'd22};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd237, 8'd145, 8'd22};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd247, 8'd151, 8'd15};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd244, 8'd145, 8'd15};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd240, 8'd137, 8'd19};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd233, 8'd127, 8'd25};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd219, 8'd113, 8'd25};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd196, 8'd94, 8'd19};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd170, 8'd72, 8'd7};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd151, 8'd57, 8'd0};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd140, 8'd21, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd118, 8'd24, 8'd0};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd111, 8'd51, 8'd25};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd127, 8'd83, 8'd58};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd128, 8'd81, 8'd53};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd130, 8'd68, 8'd29};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd162, 8'd93, 8'd36};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd206, 8'd138, 8'd67};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd209, 8'd144, 8'd54};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd220, 8'd157, 8'd64};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd225, 8'd162, 8'd65};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd218, 8'd154, 8'd56};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd208, 8'd139, 8'd44};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd203, 8'd127, 8'd41};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd196, 8'd113, 8'd35};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd189, 8'd101, 8'd29};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd178, 8'd99, 8'd43};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd176, 8'd99, 8'd45};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd169, 8'd96, 8'd45};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd148, 8'd84, 8'd40};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd144, 8'd90, 8'd56};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd156, 8'd114, 8'd90};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd210, 8'd178, 8'd163};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd217, 8'd193, 8'd183};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd240, 8'd225, 8'd206};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd244, 8'd241, 8'd236};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd210, 8'd218, 8'd229};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd187, 8'd199, 8'd213};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd198, 8'd202, 8'd211};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd238, 8'd240, 8'd239};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd244, 8'd250, 8'd248};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd216, 8'd230, 8'd230};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd213, 8'd209, 8'd210};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd205, 8'd201, 8'd198};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd176, 8'd169, 8'd163};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd149, 8'd133, 8'd120};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd140, 8'd107, 8'd88};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd130, 8'd74, 8'd47};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd123, 8'd48, 8'd16};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd133, 8'd45, 8'd9};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd158, 8'd64, 8'd28};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd145, 8'd52, 8'd19};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd121, 8'd32, 8'd0};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd123, 8'd34, 8'd4};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd149, 8'd58, 8'd27};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd163, 8'd66, 8'd31};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd158, 8'd56, 8'd16};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd156, 8'd50, 8'd8};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd168, 8'd64, 8'd25};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd148, 8'd55, 8'd12};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd193, 8'd106, 8'd61};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd162, 8'd71, 8'd26};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd169, 8'd66, 8'd25};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd171, 8'd62, 8'd21};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd155, 8'd54, 8'd10};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd146, 8'd55, 8'd8};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd146, 8'd55, 8'd8};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd138, 8'd49, 8'd7};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd128, 8'd39, 8'd9};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd119, 8'd33, 8'd10};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd121, 8'd39, 8'd18};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd128, 8'd52, 8'd28};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd128, 8'd59, 8'd26};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd123, 8'd57, 8'd22};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd133, 8'd96, 8'd78};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd142, 8'd118, 8'd106};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd154, 8'd146, 8'd143};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd156, 8'd165, 8'd170};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd153, 8'd171, 8'd181};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd149, 8'd167, 8'd179};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd146, 8'd159, 8'd168};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd144, 8'd151, 8'd161};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd147, 8'd163, 8'd179};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd141, 8'd158, 8'd174};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd149, 8'd167, 8'd179};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd142, 8'd157, 8'd162};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd156, 8'd161, 8'd155};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd169, 8'd158, 8'd138};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd172, 8'd146, 8'd113};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd158, 8'd123, 8'd83};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd166, 8'd103, 8'd49};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd161, 8'd90, 8'd36};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd154, 8'd73, 8'd20};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd156, 8'd65, 8'd12};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd162, 8'd69, 8'd12};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd166, 8'd77, 8'd17};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd165, 8'd84, 8'd19};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd161, 8'd86, 8'd18};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd186, 8'd103, 8'd35};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd173, 8'd99, 8'd28};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd168, 8'd102, 8'd26};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd172, 8'd104, 8'd31};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd169, 8'd94, 8'd29};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd151, 8'd78, 8'd25};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd135, 8'd77, 8'd31};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd130, 8'd86, 8'd41};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd124, 8'd81, 8'd46};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd115, 8'd61, 8'd27};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd116, 8'd41, 8'd9};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd134, 8'd40, 8'd2};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd161, 8'd57, 8'd6};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd186, 8'd79, 8'd7};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd204, 8'd103, 8'd11};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd216, 8'd119, 8'd14};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd236, 8'd128, 8'd20};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd245, 8'd140, 8'd23};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd250, 8'd146, 8'd23};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd245, 8'd143, 8'd15};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd239, 8'd136, 8'd17};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd230, 8'd127, 8'd24};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd215, 8'd111, 8'd26};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd201, 8'd95, 8'd21};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd205, 8'd68, 8'd32};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd189, 8'd44, 8'd15};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd189, 8'd32, 8'd17};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd192, 8'd23, 8'd28};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd184, 8'd17, 8'd27};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd172, 8'd19, 8'd11};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd160, 8'd27, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd238, 8'd118, 8'd42};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd249, 8'd163, 8'd62};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd242, 8'd165, 8'd27};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd192, 8'd108, 8'd18};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd96, 8'd1, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd114, 8'd19, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd134, 8'd37, 8'd5};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd148, 8'd49, 8'd17};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd162, 8'd66, 8'd8};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd191, 8'd89, 8'd14};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd199, 8'd96, 8'd21};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd209, 8'd106, 8'd29};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd217, 8'd111, 8'd33};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd220, 8'd114, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd224, 8'd116, 8'd28};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd230, 8'd121, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd235, 8'd126, 8'd33};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd235, 8'd121, 8'd24};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd234, 8'd120, 8'd23};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd232, 8'd120, 8'd20};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd231, 8'd118, 8'd16};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd234, 8'd117, 8'd14};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd238, 8'd115, 8'd12};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd244, 8'd112, 8'd12};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd248, 8'd112, 8'd12};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd244, 8'd123, 8'd8};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd253, 8'd129, 8'd17};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd133, 8'd22};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd134, 8'd20};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd252, 8'd133, 8'd13};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd247, 8'd140, 8'd10};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd153, 8'd12};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd254, 8'd164, 8'd16};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd247, 8'd160, 8'd18};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd251, 8'd170, 8'd37};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd243, 8'd175, 8'd64};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd98};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd243, 8'd210, 8'd156};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd218};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd79: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd182};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd246, 8'd208, 8'd137};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd236, 8'd183, 8'd71};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd236, 8'd164, 8'd17};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd246, 8'd159, 8'd0};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd0};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd13};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd25};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd29};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd253, 8'd147, 8'd25};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd253, 8'd138, 8'd21};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd130, 8'd20};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd126, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd122, 8'd25};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd116, 8'd25};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd111, 8'd21};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd117, 8'd21};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd250, 8'd110, 8'd15};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd236, 8'd98, 8'd7};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd220, 8'd89, 8'd0};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd210, 8'd86, 8'd0};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd208, 8'd89, 8'd5};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd211, 8'd96, 8'd15};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd214, 8'd101, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd205, 8'd109, 8'd23};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd201, 8'd106, 8'd22};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd195, 8'd99, 8'd22};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd184, 8'd90, 8'd20};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd170, 8'd73, 8'd18};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd155, 8'd58, 8'd16};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd141, 8'd43, 8'd14};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd134, 8'd35, 8'd14};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd113, 8'd0, 8'd18};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd160, 8'd71, 8'd15};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd226, 8'd164, 8'd29};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd220, 8'd164, 8'd17};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd222, 8'd142, 8'd47};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd174, 8'd51, 8'd18};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd190, 8'd27, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd212, 8'd25, 8'd20};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd181, 8'd19, 8'd16};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd188, 8'd36, 8'd13};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd201, 8'd65, 8'd15};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd212, 8'd96, 8'd13};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd222, 8'd119, 8'd14};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd227, 8'd134, 8'd13};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd228, 8'd140, 8'd14};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd226, 8'd141, 8'd14};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd16};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd19};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd254, 8'd138, 8'd25};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd248, 8'd130, 8'd32};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd235, 8'd119, 8'd34};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd213, 8'd99, 8'd28};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd187, 8'd77, 8'd16};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd168, 8'd62, 8'd4};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd173, 8'd43, 8'd9};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd129, 8'd29, 8'd0};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd106, 8'd41, 8'd13};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd121, 8'd75, 8'd51};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd129, 8'd82, 8'd56};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd121, 8'd63, 8'd26};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd133, 8'd68, 8'd14};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd162, 8'd94, 8'd29};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd194, 8'd118, 8'd56};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd204, 8'd134, 8'd65};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd209, 8'd143, 8'd67};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd200, 8'd137, 8'd57};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd189, 8'd128, 8'd47};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd183, 8'd119, 8'd45};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd176, 8'd107, 8'd40};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd167, 8'd96, 8'd34};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd170, 8'd98, 8'd50};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd172, 8'd104, 8'd57};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd184, 8'd121, 8'd80};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd196, 8'd143, 8'd109};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd214, 8'd176, 8'd153};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd216, 8'd194, 8'd181};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd227, 8'd217, 8'd215};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd197, 8'd195, 8'd200};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd216, 8'd214, 8'd202};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd206, 8'd214, 8'd216};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd192, 8'd210, 8'd224};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd229, 8'd245, 8'd255};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd226, 8'd233, 8'd241};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd231, 8'd233, 8'd230};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd223, 8'd233, 8'd225};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd195, 8'd212, 8'd206};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd190, 8'd171, 8'd175};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd181, 8'd163, 8'd163};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd147, 8'd123, 8'd119};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd118, 8'd84, 8'd72};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd121, 8'd66, 8'd45};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd131, 8'd52, 8'd21};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd151, 8'd49, 8'd9};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd182, 8'd65, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd175, 8'd69, 8'd29};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd159, 8'd61, 8'd24};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd132, 8'd42, 8'd15};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd126, 8'd44, 8'd20};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd148, 8'd64, 8'd40};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd159, 8'd68, 8'd39};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd157, 8'd55, 8'd17};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd159, 8'd50, 8'd7};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd171, 8'd65, 8'd23};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd150, 8'd55, 8'd9};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd192, 8'd106, 8'd57};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd161, 8'd70, 8'd23};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd168, 8'd67, 8'd25};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd170, 8'd64, 8'd24};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd12};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd142, 8'd56, 8'd9};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd137, 8'd55, 8'd8};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd138, 8'd53, 8'd14};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd129, 8'd40, 8'd10};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd117, 8'd25, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd120, 8'd28, 8'd3};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd136, 8'd47, 8'd17};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd145, 8'd60, 8'd21};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd144, 8'd60, 8'd14};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd123, 8'd65, 8'd43};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd116, 8'd70, 8'd55};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd121, 8'd96, 8'd92};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd144, 8'd139, 8'd145};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd163, 8'd169, 8'd181};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd166, 8'd173, 8'd189};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd163, 8'd165, 8'd180};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd163, 8'd159, 8'd173};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd144, 8'd141, 8'd160};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd149, 8'd154, 8'd176};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd132, 8'd148, 8'd173};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd126, 8'd152, 8'd177};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd124, 8'd151, 8'd170};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd139, 8'd157, 8'd167};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd169, 8'd178, 8'd177};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd154, 8'd155, 8'd147};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd190, 8'd142, 8'd93};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd180, 8'd124, 8'd75};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd166, 8'd98, 8'd51};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd159, 8'd82, 8'd36};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd157, 8'd79, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd155, 8'd82, 8'd29};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd149, 8'd84, 8'd26};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd143, 8'd85, 8'd22};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd175, 8'd86, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd163, 8'd83, 8'd22};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd160, 8'd86, 8'd23};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd164, 8'd88, 8'd26};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd159, 8'd76, 8'd22};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd143, 8'd62, 8'd15};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd136, 8'd69, 8'd27};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd140, 8'd87, 8'd47};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd120, 8'd81, 8'd40};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd109, 8'd55, 8'd17};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd112, 8'd37, 8'd0};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd140, 8'd43, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd170, 8'd63, 8'd7};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd191, 8'd83, 8'd8};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd208, 8'd105, 8'd12};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd221, 8'd124, 8'd17};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd243, 8'd126, 8'd13};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd252, 8'd136, 8'd17};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd255, 8'd141, 8'd14};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd249, 8'd136, 8'd6};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd239, 8'd126, 8'd4};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd230, 8'd114, 8'd11};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd213, 8'd97, 8'd14};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd197, 8'd79, 8'd9};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd185, 8'd39, 8'd24};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd176, 8'd22, 8'd10};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd187, 8'd22, 8'd16};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd195, 8'd22, 8'd28};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd184, 8'd17, 8'd25};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd168, 8'd17, 8'd6};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd154, 8'd26, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd237, 8'd125, 8'd49};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd251, 8'd162, 8'd70};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd240, 8'd159, 8'd28};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd195, 8'd107, 8'd18};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd108, 8'd12, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd124, 8'd28, 8'd4};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd130, 8'd33, 8'd1};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd142, 8'd43, 8'd12};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd164, 8'd67, 8'd16};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd185, 8'd72, 8'd2};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd193, 8'd79, 8'd9};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd203, 8'd85, 8'd15};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd207, 8'd86, 8'd15};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd208, 8'd84, 8'd10};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd210, 8'd83, 8'd4};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd215, 8'd84, 8'd2};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd218, 8'd88, 8'd2};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd241, 8'd90, 8'd7};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd244, 8'd96, 8'd10};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd106, 8'd14};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd251, 8'd117, 8'd20};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd124, 8'd20};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd127, 8'd21};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd127, 8'd19};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd127, 8'd16};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd246, 8'd148, 8'd13};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd246, 8'd145, 8'd13};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd249, 8'd144, 8'd16};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd253, 8'd148, 8'd21};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd27};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd24};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd20};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd243, 8'd165, 8'd13};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd17};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd250, 8'd163, 8'd50};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd249, 8'd191, 8'd117};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd192};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd80: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd244, 8'd217, 8'd170};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd235, 8'd196, 8'd103};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd233, 8'd179, 8'd47};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd242, 8'd167, 8'd14};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd0};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd0};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd254, 8'd152, 8'd24};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd253, 8'd151, 8'd25};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd252, 8'd150, 8'd24};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd250, 8'd148, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd248, 8'd145, 8'd24};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd246, 8'd143, 8'd24};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd243, 8'd142, 8'd24};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd242, 8'd141, 8'd25};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd118, 8'd25};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd119, 8'd28};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd117, 8'd28};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd252, 8'd114, 8'd25};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd238, 8'd104, 8'd15};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd222, 8'd92, 8'd6};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd206, 8'd80, 8'd0};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd196, 8'd72, 8'd0};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd197, 8'd64, 8'd0};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd197, 8'd63, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd195, 8'd62, 8'd0};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd188, 8'd57, 8'd1};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd176, 8'd49, 8'd8};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd157, 8'd37, 8'd10};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd140, 8'd27, 8'd11};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd129, 8'd21, 8'd11};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd115, 8'd25, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd149, 8'd54, 8'd6};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd245, 8'd156, 8'd54};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd249, 8'd164, 8'd21};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd238, 8'd147, 8'd33};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd171, 8'd52, 8'd12};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd173, 8'd17, 8'd21};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd203, 8'd25, 8'd25};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd202, 8'd33, 8'd38};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd188, 8'd26, 8'd23};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd180, 8'd30, 8'd13};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd188, 8'd57, 8'd15};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd199, 8'd84, 8'd17};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd206, 8'd108, 8'd11};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd214, 8'd128, 8'd9};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd225, 8'd144, 8'd13};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd244, 8'd141, 8'd23};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd248, 8'd142, 8'd20};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd246, 8'd137, 8'd10};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd238, 8'd126, 8'd0};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd232, 8'd119, 8'd1};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd223, 8'd109, 8'd12};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd206, 8'd90, 8'd13};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd185, 8'd71, 8'd8};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd160, 8'd44, 8'd5};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd136, 8'd32, 8'd0};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd117, 8'd33, 8'd0};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd120, 8'd51, 8'd18};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd130, 8'd71, 8'd39};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd137, 8'd78, 8'd44};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd141, 8'd77, 8'd41};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd144, 8'd76, 8'd39};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd166, 8'd103, 8'd62};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd180, 8'd104, 8'd52};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd185, 8'd100, 8'd36};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd188, 8'd107, 8'd44};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd173, 8'd103, 8'd51};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd156, 8'd98, 8'd58};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd146, 8'd92, 8'd56};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd158, 8'd102, 8'd65};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd145, 8'd110, 8'd68};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd170, 8'd141, 8'd107};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd196, 8'd178, 8'd154};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd220, 8'd216, 8'd204};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd222, 8'd228, 8'd226};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd213, 8'd228, 8'd233};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd207, 8'd225, 8'd237};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd177, 8'd196, 8'd210};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd194, 8'd214, 8'd212};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd212, 8'd232, 8'd231};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd214, 8'd232, 8'd236};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd226, 8'd241, 8'd246};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd222, 8'd232, 8'd234};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd212, 8'd217, 8'd213};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd182, 8'd182, 8'd172};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd178, 8'd176, 8'd161};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd158, 8'd121, 8'd102};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd132, 8'd89, 8'd57};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd123, 8'd69, 8'd23};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd129, 8'd61, 8'd14};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd148, 8'd64, 8'd27};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd152, 8'd58, 8'd24};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd154, 8'd57, 8'd14};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd192, 8'd92, 8'd40};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd173, 8'd70, 8'd25};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd166, 8'd74, 8'd37};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd127, 8'd43, 8'd15};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd122, 8'd37, 8'd6};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd166, 8'd70, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd178, 8'd75, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd146, 8'd45, 8'd3};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd157, 8'd61, 8'd23};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd161, 8'd62, 8'd23};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd164, 8'd65, 8'd26};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd189, 8'd90, 8'd49};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd175, 8'd76, 8'd35};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd177, 8'd78, 8'd36};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd165, 8'd66, 8'd24};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd152, 8'd54, 8'd9};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd158, 8'd60, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd157, 8'd59, 8'd14};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd158, 8'd62, 8'd24};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd137, 8'd48, 8'd18};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd114, 8'd28, 8'd3};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd120, 8'd32, 8'd8};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd145, 8'd52, 8'd19};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd158, 8'd59, 8'd17};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd162, 8'd57, 8'd9};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd133, 8'd52, 8'd5};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd125, 8'd55, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd111, 8'd53, 8'd29};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd119, 8'd72, 8'd54};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd150, 8'd113, 8'd97};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd165, 8'd146, 8'd139};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd159, 8'd168, 8'd175};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd156, 8'd187, 8'd207};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd150, 8'd163, 8'd182};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd147, 8'd162, 8'd185};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd138, 8'd156, 8'd180};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd147, 8'd169, 8'd193};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd143, 8'd168, 8'd188};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd129, 8'd156, 8'd167};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd136, 8'd164, 8'd165};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd142, 8'd168, 8'd165};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd155, 8'd166, 8'd158};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd168, 8'd169, 8'd163};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd181, 8'd166, 8'd159};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd166, 8'd134, 8'd121};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd151, 8'd101, 8'd74};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd137, 8'd75, 8'd28};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd150, 8'd81, 8'd16};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd163, 8'd90, 8'd13};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd134, 8'd62, 8'd14};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd144, 8'd55, 8'd13};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd159, 8'd55, 8'd18};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd150, 8'd48, 8'd10};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd143, 8'd59, 8'd22};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd130, 8'd65, 8'd27};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd141, 8'd85, 8'd52};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd132, 8'd77, 8'd47};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd116, 8'd52, 8'd14};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd121, 8'd50, 8'd6};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd132, 8'd49, 8'd0};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd150, 8'd55, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd174, 8'd70, 8'd0};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd198, 8'd91, 8'd0};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd219, 8'd113, 8'd3};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd231, 8'd126, 8'd9};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd224, 8'd135, 8'd9};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd226, 8'd141, 8'd16};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd221, 8'd137, 8'd15};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd206, 8'd120, 8'd9};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd199, 8'd102, 8'd8};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd199, 8'd86, 8'd16};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd196, 8'd66, 8'd17};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd187, 8'd47, 8'd12};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd201, 8'd36, 8'd34};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd187, 8'd33, 8'd25};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd174, 8'd25, 8'd19};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd164, 8'd11, 8'd16};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd167, 8'd10, 8'd21};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd170, 8'd16, 8'd14};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd161, 8'd28, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd250, 8'd136, 8'd73};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd254, 8'd160, 8'd36};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd247, 8'd159, 8'd36};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd188, 8'd98, 8'd36};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd107, 8'd16, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd108, 8'd17, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd127, 8'd26, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd149, 8'd39, 8'd6};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd160, 8'd48, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd202, 8'd39, 8'd8};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd208, 8'd45, 8'd12};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd214, 8'd55, 8'd15};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd219, 8'd61, 8'd14};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd222, 8'd65, 8'd10};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd229, 8'd73, 8'd12};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd237, 8'd84, 8'd16};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd245, 8'd92, 8'd22};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd121, 8'd6};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd125, 8'd8};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd131, 8'd12};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd138, 8'd16};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd143, 8'd21};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd252, 8'd148, 8'd23};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd249, 8'd151, 8'd24};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd247, 8'd153, 8'd27};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd242, 8'd165, 8'd37};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd248, 8'd162, 8'd25};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd11};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd1};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd3};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd245, 8'd163, 8'd19};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd232, 8'd170, 8'd37};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd223, 8'd173, 8'd50};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd233, 8'd213, 8'd150};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd237, 8'd221, 8'd169};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd240, 8'd235, 8'd197};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd81: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd200};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd156};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd249, 8'd195, 8'd107};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd237, 8'd170, 8'd63};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd230, 8'd155, 8'd38};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd16};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd18};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd21};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd24};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd27};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd27};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd253, 8'd144, 8'd27};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd250, 8'd140, 8'd25};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd240, 8'd148, 8'd11};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd242, 8'd148, 8'd16};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd248, 8'd146, 8'd22};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd251, 8'd139, 8'd27};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd251, 8'd127, 8'd27};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd245, 8'd114, 8'd24};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd241, 8'd102, 8'd21};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd236, 8'd93, 8'd15};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd220, 8'd75, 8'd0};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd218, 8'd72, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd214, 8'd68, 8'd0};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd202, 8'd59, 8'd0};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd185, 8'd48, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd165, 8'd37, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd148, 8'd25, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd137, 8'd19, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd114, 8'd22, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd145, 8'd50, 8'd2};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd246, 8'd154, 8'd51};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd240, 8'd149, 8'd34};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd173, 8'd54, 8'd14};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd170, 8'd16, 8'd18};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd198, 8'd20, 8'd20};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd186, 8'd23, 8'd26};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd191, 8'd32, 8'd29};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd189, 8'd35, 8'd23};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd184, 8'd41, 8'd11};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd188, 8'd61, 8'd8};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd206, 8'd96, 8'd17};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd218, 8'd124, 8'd24};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd220, 8'd136, 8'd22};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd232, 8'd142, 8'd22};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd236, 8'd148, 8'd22};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd233, 8'd149, 8'd15};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd226, 8'd144, 8'd8};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd221, 8'd136, 8'd9};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd215, 8'd124, 8'd17};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd198, 8'd100, 8'd13};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd179, 8'd77, 8'd3};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd169, 8'd61, 8'd22};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd145, 8'd49, 8'd9};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd124, 8'd44, 8'd7};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd122, 8'd58, 8'd23};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd130, 8'd74, 8'd41};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd134, 8'd80, 8'd46};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd139, 8'd80, 8'd46};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd144, 8'd81, 8'd46};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd138, 8'd74, 8'd36};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd160, 8'd86, 8'd37};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd167, 8'd87, 8'd28};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd161, 8'd84, 8'd28};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd147, 8'd88, 8'd44};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd148, 8'd103, 8'd72};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd127, 8'd101};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd199, 8'd158, 8'd130};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd208, 8'd195, 8'd176};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd218, 8'd209, 8'd194};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd213, 8'd210, 8'd201};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd213, 8'd218, 8'd212};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd210, 8'd219, 8'd218};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd210, 8'd220, 8'd222};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd216, 8'd226, 8'd228};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd201, 8'd211, 8'd212};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd202, 8'd222, 8'd220};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd212, 8'd228, 8'd227};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd218};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd215, 8'd220, 8'd224};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd210, 8'd208, 8'd209};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd192, 8'd183, 8'd178};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd145, 8'd128, 8'd118};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd124, 8'd105, 8'd90};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd146, 8'd90, 8'd75};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd138, 8'd79, 8'd49};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd148, 8'd79, 8'd37};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd163, 8'd80, 8'd38};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd178, 8'd84, 8'd50};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd172, 8'd69, 8'd38};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd155, 8'd49, 8'd9};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd171, 8'd65, 8'd15};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd177, 8'd72, 8'd27};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd166, 8'd72, 8'd36};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd130, 8'd46, 8'd18};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd124, 8'd37, 8'd7};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd169, 8'd71, 8'd32};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd182, 8'd77, 8'd32};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd149, 8'd48, 8'd6};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd159, 8'd63, 8'd25};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd165, 8'd63, 8'd25};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd165, 8'd63, 8'd25};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd188, 8'd86, 8'd46};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd173, 8'd71, 8'd31};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd175, 8'd74, 8'd32};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd165, 8'd64, 8'd22};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd156, 8'd55, 8'd11};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd160, 8'd59, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd160, 8'd59, 8'd13};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd159, 8'd63, 8'd23};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd140, 8'd49, 8'd20};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd116, 8'd30, 8'd5};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd119, 8'd31, 8'd7};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd144, 8'd51, 8'd20};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd159, 8'd60, 8'd19};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd160, 8'd58, 8'd9};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd145, 8'd51, 8'd0};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd142, 8'd59, 8'd17};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd126, 8'd53, 8'd21};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd114, 8'd49, 8'd21};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd123, 8'd63, 8'd37};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd129, 8'd86, 8'd67};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd138, 8'd121, 8'd113};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd153, 8'd157, 8'd160};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd166, 8'd183, 8'd190};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd167, 8'd185, 8'd195};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd156, 8'd174, 8'd188};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd154, 8'd173, 8'd190};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd143, 8'd162, 8'd179};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd129, 8'd148, 8'd163};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd140, 8'd160, 8'd169};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd144, 8'd163, 8'd169};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd139, 8'd158, 8'd162};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd151, 8'd162, 8'd168};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd171, 8'd168, 8'd175};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd187, 8'd168, 8'd170};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd194, 8'd161, 8'd152};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd178, 8'd132, 8'd108};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd154, 8'd101, 8'd61};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd132, 8'd74, 8'd24};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd127, 8'd57, 8'd8};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd134, 8'd50, 8'd6};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd150, 8'd51, 8'd12};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd142, 8'd46, 8'd8};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd142, 8'd64, 8'd25};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd136, 8'd76, 8'd39};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd140, 8'd87, 8'd55};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd119, 8'd65, 8'd37};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd114, 8'd46, 8'd9};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd121, 8'd48, 8'd5};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd136, 8'd55, 8'd0};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd155, 8'd68, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd178, 8'd86, 8'd1};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd200, 8'd108, 8'd9};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd219, 8'd129, 8'd19};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd227, 8'd140, 8'd25};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd228, 8'd151, 8'd33};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd223, 8'd146, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd223, 8'd143, 8'd32};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd221, 8'd133, 8'd35};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd209, 8'd106, 8'd27};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd194, 8'd71, 8'd14};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd188, 8'd48, 8'd12};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd193, 8'd43, 8'd19};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd195, 8'd31, 8'd32};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd182, 8'd29, 8'd24};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd169, 8'd21, 8'd17};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd160, 8'd9, 8'd14};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd165, 8'd8, 8'd19};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd167, 8'd15, 8'd10};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd163, 8'd31, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd249, 8'd136, 8'd66};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd245, 8'd154, 8'd22};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd237, 8'd152, 8'd23};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd181, 8'd91, 8'd28};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd106, 8'd13, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd111, 8'd15, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd130, 8'd24, 8'd10};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd155, 8'd37, 8'd27};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd169, 8'd49, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd187, 8'd60, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd195, 8'd68, 8'd0};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd205, 8'd79, 8'd3};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd213, 8'd88, 8'd4};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd221, 8'd96, 8'd4};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd229, 8'd105, 8'd7};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd240, 8'd117, 8'd13};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd249, 8'd127, 8'd18};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd250, 8'd128, 8'd19};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd133, 8'd22};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd28};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd146, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd26};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd254, 8'd146, 8'd20};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd249, 8'd144, 8'd17};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd252, 8'd170, 8'd8};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd248, 8'd164, 8'd4};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd6};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd237, 8'd153, 8'd18};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd235, 8'd162, 8'd49};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd236, 8'd179, 8'd90};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd241, 8'd198, 8'd130};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd243, 8'd210, 8'd157};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd82: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd254, 8'd231, 8'd215};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd245, 8'd213, 8'd174};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd238, 8'd203, 8'd149};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd224, 8'd156, 8'd31};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd229, 8'd158, 8'd32};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd240, 8'd163, 8'd35};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd248, 8'd165, 8'd33};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd29};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd22};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd15};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd9};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd237, 8'd166, 8'd0};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd241, 8'd165, 8'd1};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd245, 8'd162, 8'd8};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd248, 8'd155, 8'd15};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd249, 8'd144, 8'd19};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd247, 8'd131, 8'd20};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd242, 8'd118, 8'd18};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd240, 8'd111, 8'd17};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd239, 8'd105, 8'd18};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd234, 8'd100, 8'd15};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd223, 8'd91, 8'd9};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd209, 8'd77, 8'd5};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd188, 8'd63, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd168, 8'd48, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd148, 8'd37, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd138, 8'd30, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd112, 8'd21, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd141, 8'd45, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd245, 8'd153, 8'd50};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd165, 8'd22};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd243, 8'd152, 8'd37};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd178, 8'd59, 8'd17};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd165, 8'd12, 8'd14};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd189, 8'd14, 8'd11};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd171, 8'd17, 8'd19};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd184, 8'd26, 8'd27};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd191, 8'd29, 8'd26};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd188, 8'd28, 8'd16};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd188, 8'd40, 8'd10};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd199, 8'd73, 8'd22};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd210, 8'd106, 8'd35};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd214, 8'd123, 8'd40};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd232, 8'd159, 8'd46};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd237, 8'd172, 8'd52};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd237, 8'd184, 8'd52};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd231, 8'd188, 8'd50};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd231, 8'd184, 8'd54};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd227, 8'd170, 8'd55};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd215, 8'd140, 8'd47};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd199, 8'd112, 8'd33};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd182, 8'd90, 8'd43};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd157, 8'd73, 8'd29};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd134, 8'd61, 8'd20};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd129, 8'd67, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd131, 8'd77, 8'd43};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd132, 8'd82, 8'd49};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd138, 8'd85, 8'd53};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd144, 8'd89, 8'd58};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd140, 8'd80, 8'd43};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd151, 8'd83, 8'd38};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd149, 8'd76, 8'd25};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd146, 8'd82, 8'd38};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd159, 8'd114, 8'd83};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd170, 8'd143, 8'd126};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd189, 8'd171, 8'd159};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd216, 8'd198, 8'd184};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd198, 8'd205, 8'd211};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd209, 8'd218, 8'd223};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd213};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd193, 8'd206, 8'd212};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd217};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd209, 8'd218, 8'd217};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd225, 8'd230, 8'd224};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd224, 8'd225, 8'd217};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd202, 8'd217, 8'd212};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd219};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd201, 8'd201, 8'd199};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd199, 8'd187, 8'd187};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd182, 8'd158, 8'd154};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd159, 8'd126, 8'd117};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd117, 8'd78, 8'd63};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd105, 8'd62, 8'd43};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd155, 8'd79, 8'd65};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd158, 8'd78, 8'd51};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd169, 8'd81, 8'd41};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd173, 8'd77, 8'd35};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd186, 8'd81, 8'd49};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd185, 8'd76, 8'd47};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd162, 8'd54, 8'd16};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd166, 8'd60, 8'd12};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd180, 8'd75, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd163, 8'd69, 8'd33};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd136, 8'd50, 8'd23};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd126, 8'd39, 8'd9};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd171, 8'd73, 8'd34};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd185, 8'd80, 8'd35};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd155, 8'd52, 8'd11};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd163, 8'd65, 8'd28};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd169, 8'd67, 8'd29};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd165, 8'd63, 8'd25};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd182, 8'd80, 8'd40};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd169, 8'd67, 8'd27};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd170, 8'd69, 8'd27};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd162, 8'd61, 8'd19};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd159, 8'd58, 8'd14};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd159, 8'd58, 8'd14};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd163, 8'd61, 8'd13};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd161, 8'd64, 8'd22};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd143, 8'd52, 8'd21};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd119, 8'd33, 8'd8};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd117, 8'd31, 8'd6};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd140, 8'd49, 8'd18};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd159, 8'd62, 8'd20};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd160, 8'd58, 8'd10};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd147, 8'd42, 8'd0};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd153, 8'd55, 8'd8};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd144, 8'd55, 8'd15};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd133, 8'd45, 8'd7};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd129, 8'd44, 8'd5};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd119, 8'd46, 8'd11};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd111, 8'd61, 8'd36};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd118, 8'd86, 8'd71};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd130, 8'd136, 8'd124};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd161, 8'd168, 8'd160};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd176, 8'd185, 8'd184};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd181, 8'd190, 8'd199};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd163, 8'd175, 8'd189};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd143, 8'd159, 8'd175};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd147, 8'd164, 8'd180};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd142, 8'd161, 8'd176};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd144, 8'd173, 8'd187};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd135, 8'd158, 8'd174};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd134, 8'd149, 8'd170};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd160, 8'd162, 8'd183};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd190, 8'd182, 8'd197};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd199, 8'd180, 8'd182};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd175, 8'd151, 8'd141};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd149, 8'd120, 8'd102};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd153, 8'd87, 8'd39};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd137, 8'd59, 8'd13};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd141, 8'd52, 8'd10};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd129, 8'd46, 8'd6};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd136, 8'd69, 8'd27};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd139, 8'd87, 8'd48};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd138, 8'd89, 8'd57};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd108, 8'd57, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd129, 8'd56, 8'd21};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd139, 8'd64, 8'd22};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd157, 8'd82, 8'd25};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd181, 8'd104, 8'd32};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd203, 8'd129, 8'd42};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd221, 8'd151, 8'd53};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd234, 8'd167, 8'd62};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd68};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd234, 8'd173, 8'd67};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd225, 8'd160, 8'd58};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd221, 8'd144, 8'd52};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd217, 8'd124, 8'd47};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd205, 8'd92, 8'd34};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd193, 8'd56, 8'd20};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd190, 8'd37, 8'd19};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd199, 8'd34, 8'd28};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd184, 8'd23, 8'd31};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd173, 8'd20, 8'd23};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd158, 8'd14, 8'd14};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd157, 8'd8, 8'd14};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd161, 8'd6, 8'd14};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd165, 8'd14, 8'd5};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd168, 8'd38, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd250, 8'd139, 8'd60};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd251, 8'd163, 8'd27};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd242, 8'd158, 8'd24};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd188, 8'd96, 8'd29};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd115, 8'd17, 8'd4};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd121, 8'd20, 8'd2};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd136, 8'd25, 8'd18};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd160, 8'd37, 8'd39};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd175, 8'd51, 8'd15};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd187, 8'd89, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd195, 8'd96, 8'd2};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd205, 8'd107, 8'd6};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd213, 8'd115, 8'd8};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd218, 8'd121, 8'd6};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd226, 8'd128, 8'd5};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd234, 8'd137, 8'd7};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd242, 8'd144, 8'd11};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd27};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd22};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd253, 8'd151, 8'd17};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd251, 8'd149, 8'd15};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd252, 8'd150, 8'd14};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd16};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd19};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd22};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd242, 8'd158, 8'd10};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd239, 8'd163, 8'd25};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd238, 8'd173, 8'd55};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd239, 8'd188, 8'd97};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd242, 8'd207, 8'd143};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd248, 8'd226, 8'd187};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd83: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd193};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd168};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd246, 8'd193, 8'd125};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd231, 8'd172, 8'd80};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd227, 8'd162, 8'd44};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd23};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd252, 8'd174, 8'd12};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd12};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd7};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd10};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd14};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd17};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd17};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd250, 8'd158, 8'd15};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd244, 8'd153, 8'd13};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd239, 8'd149, 8'd11};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd237, 8'd137, 8'd26};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd231, 8'd130, 8'd24};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd220, 8'd118, 8'd20};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd202, 8'd100, 8'd16};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd183, 8'd81, 8'd15};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd161, 8'd65, 8'd17};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd144, 8'd51, 8'd18};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd133, 8'd45, 8'd21};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd117, 8'd21, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd138, 8'd40, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd245, 8'd152, 8'd48};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd249, 8'd164, 8'd19};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd247, 8'd156, 8'd39};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd184, 8'd67, 8'd24};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd160, 8'd10, 8'd9};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd182, 8'd9, 8'd5};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd162, 8'd16, 8'd16};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd165, 8'd11, 8'd13};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd179, 8'd12, 8'd19};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd196, 8'd23, 8'd27};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd198, 8'd35, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd193, 8'd51, 8'd27};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd197, 8'd78, 8'd38};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd205, 8'd104, 8'd52};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd219, 8'd149, 8'd61};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd224, 8'd170, 8'd72};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd226, 8'd193, 8'd80};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd225, 8'd206, 8'd85};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd230, 8'd211, 8'd91};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd233, 8'd199, 8'd92};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd226, 8'd169, 8'd80};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd214, 8'd143, 8'd65};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd197, 8'd116, 8'd63};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd172, 8'd96, 8'd46};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd148, 8'd77, 8'd31};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd136, 8'd75, 8'd31};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd132, 8'd76, 8'd39};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd130, 8'd80, 8'd47};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd135, 8'd86, 8'd56};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd141, 8'd94, 8'd66};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd150, 8'd94, 8'd57};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd147, 8'd82, 8'd40};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd143, 8'd76, 8'd33};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd154, 8'd100, 8'd66};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd189, 8'd157, 8'd142};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd179, 8'd171, 8'd168};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd173, 8'd174, 8'd176};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd182, 8'd186, 8'd185};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd186, 8'd194, 8'd205};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd202, 8'd212, 8'd224};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd192, 8'd206, 8'd217};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd196, 8'd210, 8'd221};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd206, 8'd221, 8'd228};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd212, 8'd223, 8'd227};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd224, 8'd230, 8'd228};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd220, 8'd225, 8'd219};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd202, 8'd205, 8'd198};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd207, 8'd202, 8'd196};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd187, 8'd170, 8'd163};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd177, 8'd144, 8'd137};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd158, 8'd111, 8'd101};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd147, 8'd89, 8'd75};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd127, 8'd62, 8'd44};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd129, 8'd63, 8'd41};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd169, 8'd83, 8'd66};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd173, 8'd86, 8'd56};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd176, 8'd83, 8'd40};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd164, 8'd65, 8'd23};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd175, 8'd72, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd184, 8'd79, 8'd49};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd168, 8'd66, 8'd28};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd169, 8'd69, 8'd20};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd183, 8'd76, 8'd32};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd160, 8'd63, 8'd28};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd142, 8'd55, 8'd28};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd128, 8'd39, 8'd9};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd174, 8'd75, 8'd36};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd189, 8'd82, 8'd38};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd162, 8'd56, 8'd16};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd165, 8'd67, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd174, 8'd70, 8'd33};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd166, 8'd62, 8'd25};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd178, 8'd74, 8'd35};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd169, 8'd65, 8'd26};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd168, 8'd65, 8'd24};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd161, 8'd58, 8'd17};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd166, 8'd63, 8'd20};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd159, 8'd56, 8'd13};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd168, 8'd63, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd163, 8'd64, 8'd22};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd150, 8'd57, 8'd24};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd125, 8'd37, 8'd13};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd115, 8'd29, 8'd4};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd137, 8'd48, 8'd18};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd160, 8'd64, 8'd24};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd157, 8'd59, 8'd14};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd150, 8'd44, 8'd0};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd8};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd148, 8'd52, 8'd14};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd14};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd160, 8'd59, 8'd17};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd142, 8'd49, 8'd8};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd106, 8'd31, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd86, 8'd28, 8'd6};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd91, 8'd63, 8'd41};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd130, 8'd103, 8'd84};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd155, 8'd135, 8'd124};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd176, 8'd165, 8'd163};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd179, 8'd180, 8'd185};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd170, 8'd184, 8'd195};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd163, 8'd189, 8'd202};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd141, 8'd173, 8'd188};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd125, 8'd159, 8'd168};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd138, 8'd172, 8'd184};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd143, 8'd171, 8'd192};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd143, 8'd167, 8'd191};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd134, 8'd150, 8'd173};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd151, 8'd160, 8'd175};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd176, 8'd179, 8'd186};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd205, 8'd205, 8'd207};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd203, 8'd142, 8'd97};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd149, 8'd78, 8'd36};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd135, 8'd58, 8'd16};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd125, 8'd54, 8'd12};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd130, 8'd76, 8'd32};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd132, 8'd87, 8'd48};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd132, 8'd83, 8'd51};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd115, 8'd59, 8'd34};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd137, 8'd57, 8'd22};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd150, 8'd73, 8'd27};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd171, 8'd99, 8'd40};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd195, 8'd129, 8'd53};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd215, 8'd155, 8'd67};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd228, 8'd175, 8'd79};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd235, 8'd187, 8'd89};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd236, 8'd192, 8'd93};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd230, 8'd179, 8'd90};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd226, 8'd163, 8'd83};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd210, 8'd130, 8'd61};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd193, 8'd89, 8'd36};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd188, 8'd61, 8'd28};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd196, 8'd49, 8'd33};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd200, 8'd36, 8'd35};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd195, 8'd24, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd172, 8'd14, 8'd28};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd162, 8'd13, 8'd19};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd149, 8'd6, 8'd8};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd153, 8'd8, 8'd15};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd157, 8'd4, 8'd9};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd162, 8'd14, 8'd0};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd173, 8'd46, 8'd0};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd252, 8'd142, 8'd57};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd25};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd233, 8'd148, 8'd19};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd181, 8'd90, 8'd20};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd116, 8'd17, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd122, 8'd22, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd137, 8'd27, 8'd4};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd162, 8'd42, 8'd25};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd178, 8'd61, 8'd7};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd197, 8'd97, 8'd3};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd206, 8'd106, 8'd8};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd218, 8'd119, 8'd17};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd229, 8'd129, 8'd18};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd235, 8'd136, 8'd19};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd243, 8'd143, 8'd19};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd252, 8'd153, 8'd24};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd29};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd253, 8'd164, 8'd0};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd4};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd12};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd253, 8'd170, 8'd16};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd247, 8'd167, 8'd20};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd239, 8'd162, 8'd20};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd229, 8'd156, 8'd17};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd224, 8'd152, 8'd14};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd244, 8'd178, 8'd100};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd246, 8'd193, 8'd125};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd251, 8'd215, 8'd163};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd254, 8'd238, 8'd202};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd84: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd217};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd186};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd247, 8'd213, 8'd142};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd231, 8'd191, 8'd95};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd215, 8'd170, 8'd55};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd205, 8'd155, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd37};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd37};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd32};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd28};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd20};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd13};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd248, 8'd161, 8'd4};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd247, 8'd160, 8'd1};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd233, 8'd154, 8'd1};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd228, 8'd146, 8'd0};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd221, 8'd132, 8'd2};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd208, 8'd113, 8'd5};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd188, 8'd92, 8'd8};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd167, 8'd71, 8'd11};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd17};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd141, 8'd45, 8'd20};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd125, 8'd27, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd138, 8'd38, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd246, 8'd150, 8'd47};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd247, 8'd163, 8'd15};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd249, 8'd160, 8'd42};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd191, 8'd76, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd159, 8'd11, 8'd7};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd177, 8'd8, 8'd1};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd155, 8'd11, 8'd10};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd155, 8'd2, 8'd5};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd167, 8'd1, 8'd11};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd188, 8'd17, 8'd26};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd200, 8'd33, 8'd40};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd196, 8'd44, 8'd39};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd191, 8'd58, 8'd41};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd191, 8'd71, 8'd46};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd203, 8'd122, 8'd67};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd210, 8'd145, 8'd79};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd214, 8'd173, 8'd91};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd217, 8'd194, 8'd100};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd227, 8'd207, 8'd110};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd236, 8'd205, 8'd114};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd235, 8'd184, 8'd105};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd225, 8'd161, 8'd90};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd203, 8'd132, 8'd70};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd182, 8'd110, 8'd51};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd159, 8'd88, 8'd34};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd146, 8'd78, 8'd29};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd136, 8'd74, 8'd33};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd130, 8'd74, 8'd41};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd131, 8'd81, 8'd54};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd138, 8'd92, 8'd68};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd142, 8'd88, 8'd52};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd132, 8'd70, 8'd33};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd134, 8'd70, 8'd34};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd150, 8'd102, 8'd79};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd190, 8'd170, 8'd163};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd155, 8'd158, 8'd165};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd131, 8'd148, 8'd156};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd140, 8'd161, 8'd166};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd187, 8'd185, 8'd188};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd202, 8'd201, 8'd206};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd197, 8'd202, 8'd208};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd200, 8'd209, 8'd218};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd203, 8'd213, 8'd222};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd204, 8'd213, 8'd220};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd210, 8'd218, 8'd221};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd200, 8'd205, 8'd208};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd195, 8'd181, 8'd168};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd190, 8'd167, 8'd153};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd161, 8'd124, 8'd108};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd157, 8'd104, 8'd88};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd156, 8'd89, 8'd72};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd159, 8'd84, 8'd63};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd139, 8'd59, 8'd36};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd138, 8'd58, 8'd33};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd164, 8'd80, 8'd54};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd173, 8'd88, 8'd49};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd177, 8'd89, 8'd39};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd165, 8'd70, 8'd22};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd173, 8'd77, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd183, 8'd86, 8'd53};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd162, 8'd69, 8'd28};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd157, 8'd67, 8'd17};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd184, 8'd77, 8'd33};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd21};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd146, 8'd59, 8'd32};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd127, 8'd36, 8'd7};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd176, 8'd74, 8'd36};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd190, 8'd81, 8'd38};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd165, 8'd59, 8'd19};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd167, 8'd67, 8'd31};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd178, 8'd74, 8'd37};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd167, 8'd63, 8'd26};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd175, 8'd71, 8'd32};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd172, 8'd68, 8'd29};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd170, 8'd67, 8'd26};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd162, 8'd59, 8'd18};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd172, 8'd69, 8'd26};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd156, 8'd53, 8'd10};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd171, 8'd65, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd166, 8'd65, 8'd21};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd155, 8'd62, 8'd29};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd130, 8'd42, 8'd18};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd113, 8'd27, 8'd4};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd135, 8'd46, 8'd16};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd160, 8'd66, 8'd28};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd156, 8'd59, 8'd16};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd14};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd146, 8'd53, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd135, 8'd44, 8'd15};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd144, 8'd47, 8'd15};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd164, 8'd62, 8'd24};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd154, 8'd56, 8'd17};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd114, 8'd33, 8'd3};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd89, 8'd23, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd115, 8'd44, 8'd16};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd123, 8'd56, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd116, 8'd59, 8'd40};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd126, 8'd86, 8'd74};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd147, 8'd130, 8'd122};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd162, 8'd168, 8'd166};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd167, 8'd195, 8'd198};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd148, 8'd187, 8'd192};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd162, 8'd189, 8'd184};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd154, 8'd184, 8'd184};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd133, 8'd166, 8'd173};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd137, 8'd171, 8'd183};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd131, 8'd163, 8'd178};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd149, 8'd177, 8'd189};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd149, 8'd172, 8'd180};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd156, 8'd175, 8'd179};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd222, 8'd168, 8'd130};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd136, 8'd74, 8'd37};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd122, 8'd57, 8'd19};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd128, 8'd69, 8'd27};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd133, 8'd86, 8'd42};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd123, 8'd78, 8'd37};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd123, 8'd69, 8'd35};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd127, 8'd60, 8'd34};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd152, 8'd67, 8'd28};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd165, 8'd85, 8'd36};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd185, 8'd114, 8'd48};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd207, 8'd146, 8'd65};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd223, 8'd169, 8'd79};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd229, 8'd182, 8'd90};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd232, 8'd186, 8'd98};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd231, 8'd186, 8'd101};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd218, 8'd158, 8'd88};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd208, 8'd137, 8'd75};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd194, 8'd99, 8'd53};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd182, 8'd63, 8'd33};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd187, 8'd47, 8'd34};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd197, 8'd42, 8'd40};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd193, 8'd29, 8'd36};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd181, 8'd14, 8'd24};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd160, 8'd8, 8'd23};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd150, 8'd7, 8'd13};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd138, 8'd2, 8'd4};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd152, 8'd9, 8'd15};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd155, 8'd4, 8'd9};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd163, 8'd16, 8'd0};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd183, 8'd56, 8'd1};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd59};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd241, 8'd155, 8'd36};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd231, 8'd145, 8'd22};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd183, 8'd90, 8'd20};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd126, 8'd27, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd136, 8'd39, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd148, 8'd46, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd173, 8'd67, 8'd19};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd193, 8'd92, 8'd2};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd224, 8'd112, 8'd4};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd233, 8'd121, 8'd11};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd243, 8'd132, 8'd17};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd249, 8'd140, 8'd23};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd251, 8'd143, 8'd19};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd252, 8'd147, 8'd19};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd21};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd23};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd29};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd247, 8'd166, 8'd25};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd228, 8'd155, 8'd24};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd214, 8'd152, 8'd33};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd214, 8'd161, 8'd55};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd228, 8'd184, 8'd89};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd245, 8'd209, 8'd123};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd144};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd85: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd235, 8'd189, 8'd114};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd235, 8'd186, 8'd107};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd237, 8'd181, 8'd94};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd239, 8'd173, 8'd77};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd241, 8'd164, 8'd58};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd40};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd243, 8'd149, 8'd25};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd243, 8'd146, 8'd16};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd244, 8'd172, 8'd10};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd244, 8'd165, 8'd10};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd239, 8'd152, 8'd11};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd231, 8'd132, 8'd12};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd215, 8'd108, 8'd10};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd193, 8'd83, 8'd6};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd174, 8'd61, 8'd5};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd163, 8'd48, 8'd3};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd136, 8'd36, 8'd10};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd141, 8'd40, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd246, 8'd151, 8'd45};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd245, 8'd159, 8'd12};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd251, 8'd162, 8'd42};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd199, 8'd84, 8'd39};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd160, 8'd15, 8'd10};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd180, 8'd13, 8'd5};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd151, 8'd3, 8'd3};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd156, 8'd6, 8'd8};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd161, 8'd4, 8'd11};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd167, 8'd7, 8'd17};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd180, 8'd23, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd197, 8'd44, 8'd46};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd196, 8'd51, 8'd46};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd186, 8'd45, 8'd35};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd195, 8'd90, 8'd60};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd201, 8'd109, 8'd68};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd205, 8'd132, 8'd77};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd209, 8'd155, 8'd85};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd220, 8'd174, 8'd96};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd232, 8'd185, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd232, 8'd176, 8'd99};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd224, 8'd162, 8'd87};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd204, 8'd134, 8'd62};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd187, 8'd114, 8'd45};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd167, 8'd92, 8'd27};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd154, 8'd77, 8'd21};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd142, 8'd68, 8'd23};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd130, 8'd64, 8'd29};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd127, 8'd71, 8'd44};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd134, 8'd84, 8'd61};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd146, 8'd92, 8'd58};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd125, 8'd65, 8'd29};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd117, 8'd54, 8'd23};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd81, 8'd63};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd187, 8'd169, 8'd169};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd154, 8'd163, 8'd172};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd129, 8'd151, 8'd162};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd131, 8'd159, 8'd163};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd197, 8'd190, 8'd184};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd202, 8'd197, 8'd193};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd204, 8'd200, 8'd199};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd205, 8'd203, 8'd206};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd192, 8'd187, 8'd191};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd186, 8'd177, 8'd178};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd187, 8'd175, 8'd175};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd162, 8'd147, 8'd144};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd167, 8'd131, 8'd109};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd173, 8'd128, 8'd105};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd160, 8'd102, 8'd78};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd165, 8'd93, 8'd68};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd163, 8'd82, 8'd55};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd158, 8'd74, 8'd48};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd132, 8'd48, 8'd22};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd127, 8'd46, 8'd19};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd163, 8'd79, 8'd45};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd173, 8'd86, 8'd41};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd177, 8'd88, 8'd32};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd165, 8'd71, 8'd19};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd174, 8'd77, 8'd35};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd182, 8'd85, 8'd52};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd160, 8'd66, 8'd28};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd155, 8'd64, 8'd17};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd184, 8'd75, 8'd32};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd145, 8'd47, 8'd12};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd149, 8'd59, 8'd33};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd123, 8'd32, 8'd3};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd174, 8'd72, 8'd34};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd189, 8'd80, 8'd37};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd167, 8'd59, 8'd20};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd168, 8'd65, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd183, 8'd76, 8'd40};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd171, 8'd64, 8'd28};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd178, 8'd72, 8'd33};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd181, 8'd75, 8'd36};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd178, 8'd72, 8'd32};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd167, 8'd61, 8'd21};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd180, 8'd74, 8'd32};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd155, 8'd49, 8'd7};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd175, 8'd68, 8'd16};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd168, 8'd65, 8'd20};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd161, 8'd67, 8'd33};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd135, 8'd48, 8'd21};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd111, 8'd25, 8'd2};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd131, 8'd44, 8'd16};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd160, 8'd68, 8'd31};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd156, 8'd60, 8'd18};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd137, 8'd49, 8'd13};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd137, 8'd52, 8'd21};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd131, 8'd45, 8'd20};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd19};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd158, 8'd58, 8'd24};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd150, 8'd52, 8'd17};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd118, 8'd34, 8'd6};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd98, 8'd30, 8'd9};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd140, 8'd45, 8'd13};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd142, 8'd51, 8'd22};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd121, 8'd40, 8'd11};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd109, 8'd43, 8'd19};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd103, 8'd58, 8'd39};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd110, 8'd93, 8'd77};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd142, 8'd145, 8'd134};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd152, 8'd169, 8'd161};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd172, 8'd178, 8'd164};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd191, 8'd202, 8'd194};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd178, 8'd200, 8'd198};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd160, 8'd189, 8'd195};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd103, 8'd136, 8'd145};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd101, 8'd134, 8'd141};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd112, 8'd141, 8'd145};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd148, 8'd174, 8'd175};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd204, 8'd157, 8'd131};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd107, 8'd53, 8'd25};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd111, 8'd55, 8'd22};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd137, 8'd85, 8'd46};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd137, 8'd94, 8'd49};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd118, 8'd69, 8'd26};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd121, 8'd53, 8'd18};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd140, 8'd54, 8'd27};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd170, 8'd79, 8'd34};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd178, 8'd96, 8'd40};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd196, 8'd122, 8'd49};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd212, 8'd148, 8'd61};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd223, 8'd164, 8'd74};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd224, 8'd168, 8'd81};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd222, 8'd165, 8'd88};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd218, 8'd159, 8'd89};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd201, 8'd120, 8'd67};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd190, 8'd95, 8'd51};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd188, 8'd70, 8'd42};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd196, 8'd58, 8'd47};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd200, 8'd48, 8'd47};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd186, 8'd30, 8'd34};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd169, 8'd14, 8'd20};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd159, 8'd8, 8'd13};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd152, 8'd4, 8'd16};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd142, 8'd3, 8'd8};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd132, 8'd0, 8'd0};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd151, 8'd12, 8'd17};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd155, 8'd6, 8'd10};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd164, 8'd18, 8'd3};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd193, 8'd66, 8'd11};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd67};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd51};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd239, 8'd153, 8'd32};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd190, 8'd96, 8'd24};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd134, 8'd36, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd140, 8'd47, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd142, 8'd52, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd163, 8'd73, 8'd13};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd185, 8'd101, 8'd2};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd219, 8'd118, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd228, 8'd129, 8'd10};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd238, 8'd142, 8'd22};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd245, 8'd152, 8'd33};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd246, 8'd157, 8'd37};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd246, 8'd162, 8'd40};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd247, 8'd167, 8'd44};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd250, 8'd172, 8'd48};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd227, 8'd164, 8'd87};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd235, 8'd175, 8'd105};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd195, 8'd135};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd168};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd200};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd86: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd247, 8'd248, 8'd214};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd248, 8'd244, 8'd207};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd247, 8'd235, 8'd193};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd247, 8'd225, 8'd176};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd246, 8'd214, 8'd157};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd247, 8'd203, 8'd140};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd248, 8'd195, 8'd127};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd248, 8'd191, 8'd120};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd219, 8'd174, 8'd73};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd222, 8'd170, 8'd71};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd222, 8'd159, 8'd64};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd215, 8'd139, 8'd53};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd199, 8'd112, 8'd35};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd175, 8'd80, 8'd14};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd152, 8'd53, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd137, 8'd36, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd147, 8'd46, 8'd18};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd145, 8'd41, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd247, 8'd150, 8'd43};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd242, 8'd156, 8'd7};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd252, 8'd164, 8'd41};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd204, 8'd92, 8'd44};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd164, 8'd20, 8'd12};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd183, 8'd19, 8'd9};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd158, 8'd4, 8'd4};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd158, 8'd8, 8'd9};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd152, 8'd8, 8'd8};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd147, 8'd4, 8'd6};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd157, 8'd14, 8'd16};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd181, 8'd33, 8'd33};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd198, 8'd44, 8'd42};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd202, 8'd45, 8'd40};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd188, 8'd56, 8'd31};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd193, 8'd68, 8'd36};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd195, 8'd84, 8'd39};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd197, 8'd101, 8'd41};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd205, 8'd123, 8'd50};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd214, 8'd143, 8'd61};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd213, 8'd147, 8'd60};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd205, 8'd141, 8'd51};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd200, 8'd129, 8'd49};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd188, 8'd110, 8'd35};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd173, 8'd89, 8'd19};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd162, 8'd73, 8'd13};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd147, 8'd61, 8'd12};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd130, 8'd54, 8'd18};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd125, 8'd61, 8'd33};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd129, 8'd72, 8'd52};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd154, 8'd100, 8'd64};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd140, 8'd77, 8'd42};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd121, 8'd58, 8'd27};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd112, 8'd65, 8'd49};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd186, 8'd166, 8'd167};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd174, 8'd181, 8'd191};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd159, 8'd182, 8'd188};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd157, 8'd183, 8'd182};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd221, 8'd227, 8'd225};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd206, 8'd210, 8'd209};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd200, 8'd199, 8'd197};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd193, 8'd182, 8'd178};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd159, 8'd136, 8'd128};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd156, 8'd118, 8'd105};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd167, 8'd119, 8'd99};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd135, 8'd79, 8'd56};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd140, 8'd83, 8'd54};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd164, 8'd99, 8'd69};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd170, 8'd95, 8'd63};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd182, 8'd98, 8'd64};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd174, 8'd85, 8'd53};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd158, 8'd71, 8'd41};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd126, 8'd45, 8'd16};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd120, 8'd44, 8'd18};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd175, 8'd81, 8'd45};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd177, 8'd82, 8'd36};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd178, 8'd79, 8'd22};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd13};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd178, 8'd68, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd185, 8'd74, 8'd46};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd168, 8'd59, 8'd26};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd23};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd183, 8'd74, 8'd31};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd138, 8'd38, 8'd4};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd150, 8'd60, 8'd34};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd122, 8'd28, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd173, 8'd69, 8'd32};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd189, 8'd78, 8'd35};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd166, 8'd58, 8'd19};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd167, 8'd64, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd184, 8'd77, 8'd41};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd172, 8'd65, 8'd29};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd180, 8'd74, 8'd35};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd189, 8'd83, 8'd44};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd185, 8'd79, 8'd39};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd172, 8'd66, 8'd26};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd186, 8'd80, 8'd38};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd152, 8'd46, 8'd4};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd179, 8'd69, 8'd16};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd171, 8'd66, 8'd21};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd167, 8'd70, 8'd37};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd138, 8'd51, 8'd24};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd109, 8'd23, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd129, 8'd42, 8'd15};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd159, 8'd69, 8'd34};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd154, 8'd61, 8'd20};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd130, 8'd41, 8'd0};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd137, 8'd51, 8'd16};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd139, 8'd52, 8'd24};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd150, 8'd55, 8'd23};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd166, 8'd62, 8'd25};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd152, 8'd50, 8'd12};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd115, 8'd28, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd95, 8'd23, 8'd1};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd125, 8'd40, 8'd1};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd146, 8'd58, 8'd20};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd147, 8'd59, 8'd21};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd137, 8'd53, 8'd19};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd105, 8'd31, 8'd2};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd85, 8'd27, 8'd5};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd113, 8'd72, 8'd54};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd138, 8'd106, 8'd93};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd159, 8'd139, 8'd130};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd181, 8'd170, 8'd164};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd171, 8'd172, 8'd174};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd157, 8'd174, 8'd181};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd98, 8'd123, 8'd130};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd100, 8'd127, 8'd134};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd111, 8'd135, 8'd139};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd148, 8'd169, 8'd172};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd194, 8'd152, 8'd138};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd99, 8'd52, 8'd34};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd116, 8'd66, 8'd41};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd139, 8'd93, 8'd57};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd133, 8'd90, 8'd45};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd115, 8'd61, 8'd15};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd124, 8'd45, 8'd6};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd155, 8'd52, 8'd21};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd164, 8'd73, 8'd20};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd171, 8'd86, 8'd22};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd184, 8'd107, 8'd27};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd194, 8'd123, 8'd33};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd199, 8'd130, 8'd39};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd197, 8'd125, 8'd43};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd192, 8'd114, 8'd48};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd187, 8'd105, 8'd49};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd190, 8'd81, 8'd42};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd193, 8'd70, 8'd39};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd203, 8'd61, 8'd47};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd210, 8'd55, 8'd53};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd199, 8'd38, 8'd44};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd171, 8'd18, 8'd23};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd150, 8'd8, 8'd7};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd142, 8'd10, 8'd5};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd146, 8'd3, 8'd9};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd137, 8'd3, 8'd2};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd127, 8'd0, 8'd0};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd152, 8'd16, 8'd18};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd155, 8'd8, 8'd14};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd165, 8'd22, 8'd8};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd203, 8'd76, 8'd25};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd75};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd251, 8'd161, 8'd39};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd234, 8'd146, 8'd20};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd185, 8'd91, 8'd17};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd132, 8'd35, 8'd2};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd137, 8'd49, 8'd1};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd137, 8'd54, 8'd12};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd156, 8'd76, 8'd41};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd178, 8'd108, 8'd36};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd201, 8'd138, 8'd58};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd213, 8'd152, 8'd72};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd228, 8'd172, 8'd95};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd239, 8'd191, 8'd115};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd244, 8'd205, 8'd130};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd143};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd252, 8'd225, 8'd154};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd162};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd87: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd182};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd240, 8'd188, 8'd148};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd215, 8'd153, 8'd112};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd186, 8'd121, 8'd81};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd169, 8'd101, 8'd62};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd154, 8'd53, 8'd25};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd148, 8'd44, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd247, 8'd150, 8'd43};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd241, 8'd155, 8'd6};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd252, 8'd164, 8'd41};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd207, 8'd95, 8'd47};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd166, 8'd23, 8'd15};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd187, 8'd23, 8'd13};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd171, 8'd13, 8'd12};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd156, 8'd6, 8'd5};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd143, 8'd5, 8'd3};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd138, 8'd9, 8'd4};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd143, 8'd11, 8'd7};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd160, 8'd17, 8'd13};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd194, 8'd36, 8'd33};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd226, 8'd58, 8'd55};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd203, 8'd55, 8'd27};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd207, 8'd63, 8'd29};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd207, 8'd70, 8'd26};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd204, 8'd81, 8'd21};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd210, 8'd104, 8'd28};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd217, 8'd129, 8'd39};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd214, 8'd142, 8'd42};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd203, 8'd140, 8'd34};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd195, 8'd123, 8'd39};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd187, 8'd106, 8'd25};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd177, 8'd86, 8'd13};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd166, 8'd71, 8'd7};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd150, 8'd56, 8'd4};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd131, 8'd47, 8'd10};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd123, 8'd54, 8'd25};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd126, 8'd65, 8'd44};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd140, 8'd86, 8'd50};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd153, 8'd90, 8'd55};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd143, 8'd80, 8'd49};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd111, 8'd62, 8'd47};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd173, 8'd152, 8'd151};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd172, 8'd177, 8'd183};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd178, 8'd197, 8'd201};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd182, 8'd207, 8'd203};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd199, 8'd222, 8'd228};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd168, 8'd183, 8'd188};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd148, 8'd152, 8'd151};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd135, 8'd120, 8'd113};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd102, 8'd65, 8'd47};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd123, 8'd63, 8'd35};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd169, 8'd89, 8'd52};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd149, 8'd58, 8'd14};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd139, 8'd71, 8'd36};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd158, 8'd82, 8'd48};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd164, 8'd79, 8'd42};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd187, 8'd95, 8'd56};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd190, 8'd98, 8'd61};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd176, 8'd90, 8'd57};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd133, 8'd56, 8'd26};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd116, 8'd46, 8'd20};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd177, 8'd74, 8'd39};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd179, 8'd74, 8'd27};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd184, 8'd75, 8'd19};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd180, 8'd64, 8'd15};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd68, 8'd34};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd193, 8'd69, 8'd45};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd173, 8'd49, 8'd23};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd175, 8'd55, 8'd21};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd183, 8'd72, 8'd29};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd134, 8'd34, 8'd0};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd150, 8'd58, 8'd33};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd119, 8'd25, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd171, 8'd67, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd188, 8'd77, 8'd34};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd167, 8'd58, 8'd19};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd165, 8'd62, 8'd27};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd185, 8'd77, 8'd41};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd174, 8'd66, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd183, 8'd75, 8'd37};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd196, 8'd88, 8'd50};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd191, 8'd83, 8'd44};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd176, 8'd68, 8'd29};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd190, 8'd83, 8'd41};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd151, 8'd44, 8'd2};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd180, 8'd70, 8'd17};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd171, 8'd66, 8'd19};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd169, 8'd72, 8'd37};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd140, 8'd53, 8'd26};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd108, 8'd24, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd127, 8'd41, 8'd14};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd160, 8'd70, 8'd36};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd154, 8'd61, 8'd20};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd147, 8'd52, 8'd4};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd148, 8'd56, 8'd15};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd145, 8'd52, 8'd18};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd155, 8'd55, 8'd19};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd173, 8'd66, 8'd24};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd159, 8'd53, 8'd11};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd118, 8'd28, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd93, 8'd17, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd111, 8'd43, 8'd0};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd130, 8'd56, 8'd9};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd144, 8'd60, 8'd16};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd156, 8'd64, 8'd23};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd135, 8'd42, 8'd8};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd104, 8'd17, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd109, 8'd31, 8'd11};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd118, 8'd44, 8'd31};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd88, 8'd50, 8'd47};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd141, 8'd112, 8'd114};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd164, 8'd153, 8'd161};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd174, 8'd178, 8'd190};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd112, 8'd128, 8'd141};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd110, 8'd128, 8'd140};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd115, 8'd132, 8'd140};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd155, 8'd170, 8'd177};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd202, 8'd165, 8'd157};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd110, 8'd68, 8'd56};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd128, 8'd82, 8'd59};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd139, 8'd96, 8'd61};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd124, 8'd81, 8'd36};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd115, 8'd54, 8'd7};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd132, 8'd43, 8'd3};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd165, 8'd52, 8'd18};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd171, 8'd76, 8'd20};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd176, 8'd87, 8'd19};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd184, 8'd103, 8'd21};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd189, 8'd114, 8'd21};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd190, 8'd115, 8'd24};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd187, 8'd104, 8'd26};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd181, 8'd88, 8'd29};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd178, 8'd77, 8'd31};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd187, 8'd58, 8'd26};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd209, 8'd69, 8'd46};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd223, 8'd66, 8'd59};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd209, 8'd43, 8'd47};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd184, 8'd19, 8'd26};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd162, 8'd12, 8'd14};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd145, 8'd13, 8'd8};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd132, 8'd14, 8'd2};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd143, 8'd3, 8'd4};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd135, 8'd3, 8'd0};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd125, 8'd0, 8'd0};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd153, 8'd19, 8'd20};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd157, 8'd10, 8'd16};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd166, 8'd22, 8'd11};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd207, 8'd81, 8'd33};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd80};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd250, 8'd162, 8'd29};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd237, 8'd149, 8'd15};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd195, 8'd101, 8'd27};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd152, 8'd57, 8'd29};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd166, 8'd80, 8'd47};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd174, 8'd93, 8'd76};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd198, 8'd123, 8'd118};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd226, 8'd161, 8'd123};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd88: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd239, 8'd222, 8'd192};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd222, 8'd191, 8'd162};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd204, 8'd157, 8'd129};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd188, 8'd126, 8'd103};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd178, 8'd107, 8'd89};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd161, 8'd61, 8'd25};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd144, 8'd46, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd242, 8'd151, 8'd37};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd235, 8'd150, 8'd21};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd254, 8'd166, 8'd56};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd220, 8'd108, 8'd45};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd176, 8'd26, 8'd12};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd195, 8'd17, 8'd33};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd158, 8'd8, 8'd7};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd152, 8'd9, 8'd5};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd142, 8'd7, 8'd1};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd139, 8'd7, 8'd2};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd142, 8'd8, 8'd5};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd155, 8'd11, 8'd11};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd169, 8'd14, 8'd20};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd179, 8'd15, 8'd24};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd199, 8'd51, 8'd49};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd199, 8'd52, 8'd45};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd197, 8'd57, 8'd42};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd195, 8'd66, 8'd37};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd196, 8'd82, 8'd32};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd198, 8'd101, 8'd32};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd201, 8'd120, 8'd31};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd204, 8'd131, 8'd29};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd210, 8'd131, 8'd36};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd203, 8'd120, 8'd28};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd190, 8'd99, 8'd16};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd175, 8'd78, 8'd7};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd160, 8'd61, 8'd2};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd147, 8'd52, 8'd8};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd139, 8'd49, 8'd15};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd135, 8'd48, 8'd21};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd148, 8'd83, 8'd53};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd139, 8'd76, 8'd41};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd127, 8'd75, 8'd38};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd130, 8'd103, 8'd74};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd175, 8'd173, 8'd161};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd167, 8'd181, 8'd181};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd169, 8'd180, 8'd182};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd190, 8'd196, 8'd196};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd208, 8'd205, 8'd224};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd158, 8'd173, 8'd180};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd154, 8'd151, 8'd146};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd125, 8'd70, 8'd50};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd141, 8'd56, 8'd19};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd145, 8'd67, 8'd18};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd170, 8'd95, 8'd53};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd150, 8'd58, 8'd33};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd158, 8'd71, 8'd28};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd156, 8'd67, 8'd23};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd152, 8'd61, 8'd17};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd163, 8'd70, 8'd26};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd187, 8'd95, 8'd54};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd98, 8'd60};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd151, 8'd67, 8'd33};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd114, 8'd33, 8'd3};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd179, 8'd80, 8'd41};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd180, 8'd77, 8'd36};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd179, 8'd72, 8'd28};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd169, 8'd58, 8'd13};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd188, 8'd75, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd190, 8'd79, 8'd36};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd162, 8'd53, 8'd14};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd174, 8'd66, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd193, 8'd70, 8'd37};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd154, 8'd45, 8'd12};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd151, 8'd58, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd126, 8'd32, 8'd4};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd159, 8'd55, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd198, 8'd85, 8'd55};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd182, 8'd70, 8'd32};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd163, 8'd58, 8'd11};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd169, 8'd66, 8'd23};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd186, 8'd80, 8'd38};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd166, 8'd57, 8'd18};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd188, 8'd78, 8'd41};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd186, 8'd76, 8'd39};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd171, 8'd64, 8'd28};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd160, 8'd61, 8'd22};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd171, 8'd73, 8'd36};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd185, 8'd75, 8'd26};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd164, 8'd57, 8'd13};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd183, 8'd81, 8'd43};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd146, 8'd51, 8'd21};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd106, 8'd15, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd138, 8'd48, 8'd22};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd160, 8'd70, 8'd43};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd161, 8'd70, 8'd41};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd142, 8'd43, 8'd4};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd143, 8'd50, 8'd16};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd41, 8'd6};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd150, 8'd61, 8'd19};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd153, 8'd57, 8'd9};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd148, 8'd53, 8'd9};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd123, 8'd38, 8'd9};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd95, 8'd22, 8'd5};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd111, 8'd37, 8'd12};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd136, 8'd52, 8'd16};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd56, 8'd12};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd157, 8'd62, 8'd18};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd134, 8'd51, 8'd11};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd115, 8'd37, 8'd1};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd134, 8'd52, 8'd12};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd149, 8'd61, 8'd15};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd114, 8'd34, 8'd0};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd112, 8'd61, 8'd40};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd162, 8'd152, 8'd150};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd161, 8'd178, 8'd186};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd128, 8'd153, 8'd160};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd134, 8'd154, 8'd161};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd142, 8'd160, 8'd170};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd159, 8'd177, 8'd191};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd188, 8'd171, 8'd145};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd113, 8'd87, 8'd60};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd123, 8'd84, 8'd53};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd135, 8'd79, 8'd44};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd138, 8'd64, 8'd25};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd129, 8'd41, 8'd1};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd142, 8'd43, 8'd1};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd177, 8'd71, 8'd29};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd176, 8'd87, 8'd29};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd174, 8'd89, 8'd24};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd181, 8'd99, 8'd25};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd194, 8'd111, 8'd31};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd198, 8'd106, 8'd33};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd191, 8'd87, 8'd26};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd191, 8'd72, 8'd29};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd198, 8'd71, 8'd38};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd223, 8'd84, 8'd79};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd209, 8'd66, 8'd62};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd190, 8'd40, 8'd39};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd176, 8'd23, 8'd25};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd167, 8'd14, 8'd16};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd156, 8'd10, 8'd11};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd144, 8'd4, 8'd3};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd134, 8'd0, 8'd0};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd143, 8'd4, 8'd9};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd148, 8'd3, 8'd0};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd146, 8'd9, 8'd0};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd152, 8'd21, 8'd11};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd174, 8'd20, 8'd28};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd198, 8'd22, 8'd25};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd225, 8'd80, 8'd35};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd67};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd233, 8'd152, 8'd17};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd228, 8'd145, 8'd41};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd183, 8'd95, 8'd31};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd141, 8'd53, 8'd13};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd143, 8'd63, 8'd26};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd164, 8'd91, 8'd50};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd192, 8'd125, 8'd83};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd228, 8'd165, 8'd124};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd229, 8'd194, 8'd166};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd89: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd252, 8'd239, 8'd161};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd249, 8'd234, 8'd153};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd240, 8'd222, 8'd138};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd227, 8'd201, 8'd116};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd209, 8'd171, 8'd88};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd190, 8'd137, 8'd59};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd174, 8'd106, 8'd35};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd163, 8'd88, 8'd21};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd161, 8'd62, 8'd23};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd144, 8'd46, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd241, 8'd151, 8'd37};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd234, 8'd151, 8'd19};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd254, 8'd168, 8'd57};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd222, 8'd110, 8'd46};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd181, 8'd31, 8'd16};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd205, 8'd24, 8'd39};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd161, 8'd9, 8'd6};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd153, 8'd8, 8'd5};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd144, 8'd7, 8'd1};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd138, 8'd6, 8'd1};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd139, 8'd7, 8'd3};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd149, 8'd9, 8'd8};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd160, 8'd11, 8'd15};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd169, 8'd12, 8'd19};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd183, 8'd33, 8'd34};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd201, 8'd53, 8'd51};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd215, 8'd73, 8'd63};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd206, 8'd74, 8'd51};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd184, 8'd67, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd175, 8'd73, 8'd11};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd185, 8'd98, 8'd18};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd202, 8'd122, 8'd33};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd196, 8'd115, 8'd23};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd195, 8'd111, 8'd21};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd191, 8'd100, 8'd17};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd179, 8'd85, 8'd13};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd163, 8'd67, 8'd6};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd148, 8'd53, 8'd5};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd137, 8'd47, 8'd10};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd132, 8'd45, 8'd15};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd127, 8'd64, 8'd33};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd134, 8'd71, 8'd36};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd127, 8'd77, 8'd40};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd123, 8'd96, 8'd69};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd163, 8'd163, 8'd153};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd169, 8'd183, 8'd184};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd177, 8'd192, 8'd197};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd194, 8'd204, 8'd205};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd229, 8'd228, 8'd246};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd169, 8'd186, 8'd193};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd149, 8'd148, 8'd143};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd119, 8'd63, 8'd46};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd136, 8'd50, 8'd15};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd143, 8'd65, 8'd16};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd169, 8'd92, 8'd50};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd144, 8'd52, 8'd27};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd159, 8'd70, 8'd28};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd156, 8'd65, 8'd21};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd151, 8'd58, 8'd14};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd163, 8'd68, 8'd24};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd184, 8'd91, 8'd50};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd96, 8'd59};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd155, 8'd69, 8'd36};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd121, 8'd38, 8'd8};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd178, 8'd79, 8'd40};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd182, 8'd79, 8'd38};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd179, 8'd72, 8'd28};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd171, 8'd60, 8'd15};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd188, 8'd75, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd189, 8'd78, 8'd35};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd163, 8'd54, 8'd15};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd175, 8'd67, 8'd31};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd193, 8'd69, 8'd35};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd157, 8'd48, 8'd15};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd152, 8'd59, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd126, 8'd32, 8'd4};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd160, 8'd56, 8'd29};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd197, 8'd84, 8'd54};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd183, 8'd71, 8'd33};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd166, 8'd59, 8'd13};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd158, 8'd55, 8'd12};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd188, 8'd81, 8'd39};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd173, 8'd64, 8'd25};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd178, 8'd66, 8'd28};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd189, 8'd79, 8'd42};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd193, 8'd86, 8'd50};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd175, 8'd73, 8'd35};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd147, 8'd49, 8'd10};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd178, 8'd75, 8'd32};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd185, 8'd86, 8'd47};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd147, 8'd52, 8'd20};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd129, 8'd39, 8'd13};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd120, 8'd34, 8'd9};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd120, 8'd32, 8'd8};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd152, 8'd61, 8'd34};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd155, 8'd62, 8'd31};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd142, 8'd43, 8'd4};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd143, 8'd50, 8'd16};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd41, 8'd6};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd150, 8'd61, 8'd21};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd11};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd148, 8'd52, 8'd10};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd123, 8'd38, 8'd9};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd95, 8'd22, 8'd5};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd111, 8'd37, 8'd12};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd137, 8'd53, 8'd17};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd56, 8'd12};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd156, 8'd61, 8'd17};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd135, 8'd50, 8'd11};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd117, 8'd37, 8'd2};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd136, 8'd53, 8'd13};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd150, 8'd59, 8'd14};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd124, 8'd44, 8'd7};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd124, 8'd73, 8'd52};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd161};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd170, 8'd187, 8'd195};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd138, 8'd163, 8'd170};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd144, 8'd164, 8'd171};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd151, 8'd169, 8'd181};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd168, 8'd185, 8'd201};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd187, 8'd166, 8'd145};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd116, 8'd88, 8'd64};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd123, 8'd82, 8'd52};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd127, 8'd68, 8'd34};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd132, 8'd57, 8'd17};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd136, 8'd47, 8'd3};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd147, 8'd49, 8'd4};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd168, 8'd65, 8'd20};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd166, 8'd76, 8'd16};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd178, 8'd89, 8'd23};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd186, 8'd98, 8'd26};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd183, 8'd92, 8'd19};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd178, 8'd79, 8'd12};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd184, 8'd72, 8'd22};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd200, 8'd76, 8'd42};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd213, 8'd81, 8'd56};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd204, 8'd65, 8'd60};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd193, 8'd50, 8'd46};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd177, 8'd29, 8'd27};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd168, 8'd15, 8'd17};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd160, 8'd10, 8'd11};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd155, 8'd9, 8'd10};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd147, 8'd7, 8'd6};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd142, 8'd4, 8'd2};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd142, 8'd1, 8'd7};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd150, 8'd2, 8'd0};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd152, 8'd10, 8'd0};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd157, 8'd24, 8'd15};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd179, 8'd24, 8'd32};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd200, 8'd24, 8'd27};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd224, 8'd82, 8'd36};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd67};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd243, 8'd162, 8'd19};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd233, 8'd147, 8'd34};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd179, 8'd91, 8'd17};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd135, 8'd48, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd138, 8'd58, 8'd9};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd152, 8'd81, 8'd25};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd167, 8'd105, 8'd44};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd194, 8'd135, 8'd75};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd209, 8'd167, 8'd83};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd229, 8'd193, 8'd109};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd246, 8'd217, 8'd137};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd250, 8'd229, 8'd150};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd247, 8'd233, 8'd158};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd250, 8'd240, 8'd169};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd254, 8'd243, 8'd177};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd254, 8'd243, 8'd179};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd90: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd244, 8'd240, 8'd192};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd243, 8'd236, 8'd158};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd248, 8'd236, 8'd152};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd254, 8'd235, 8'd166};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd188};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd204};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd252, 8'd253, 8'd211};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd253, 8'd255, 8'd215};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd220};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd253, 8'd255, 8'd224};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd223};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd251, 8'd255, 8'd218};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd250, 8'd252, 8'd212};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd248, 8'd249, 8'd207};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd217};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd215};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd211};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd204};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd197};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd253, 8'd239, 8'd190};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd253, 8'd237, 8'd186};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd253, 8'd236, 8'd184};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd253, 8'd229, 8'd155};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd251, 8'd227, 8'd153};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd248, 8'd225, 8'd149};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd246, 8'd221, 8'd141};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd242, 8'd215, 8'd134};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd238, 8'd212, 8'd128};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd236, 8'd208, 8'd124};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd234, 8'd207, 8'd120};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd241, 8'd211, 8'd87};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd239, 8'd208, 8'd83};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd235, 8'd201, 8'd77};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd227, 8'd187, 8'd65};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd215, 8'd164, 8'd49};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd201, 8'd136, 8'd32};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd189, 8'd110, 8'd17};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd181, 8'd95, 8'd8};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd168, 8'd64, 8'd25};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd148, 8'd50, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd40};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd232, 8'd156, 8'd19};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd251, 8'd171, 8'd56};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd222, 8'd115, 8'd47};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd189, 8'd38, 8'd21};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd218, 8'd33, 8'd47};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd169, 8'd11, 8'd10};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd161, 8'd9, 8'd6};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd148, 8'd6, 8'd2};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd138, 8'd5, 8'd0};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd136, 8'd4, 8'd0};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd140, 8'd6, 8'd3};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd148, 8'd8, 8'd7};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd154, 8'd10, 8'd10};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd164, 8'd14, 8'd16};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd192, 8'd43, 8'd45};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd219, 8'd74, 8'd71};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd217, 8'd79, 8'd66};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd191, 8'd66, 8'd36};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd171, 8'd60, 8'd14};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd174, 8'd76, 8'd13};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd183, 8'd95, 8'd21};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd185, 8'd99, 8'd12};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd190, 8'd101, 8'd17};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd189, 8'd98, 8'd17};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd179, 8'd87, 8'd14};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd162, 8'd68, 8'd4};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd146, 8'd55, 8'd2};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd138, 8'd49, 8'd7};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd135, 8'd50, 8'd13};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd109, 8'd48, 8'd17};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd130, 8'd70, 8'd34};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd132, 8'd82, 8'd47};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd120, 8'd92, 8'd68};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd153, 8'd153, 8'd145};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd166, 8'd181, 8'd186};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd177, 8'd196, 8'd202};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd186, 8'd200, 8'd203};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd185, 8'd187, 8'd202};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd146, 8'd164, 8'd168};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd141, 8'd140, 8'd135};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd127, 8'd71, 8'd56};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd139, 8'd53, 8'd20};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd143, 8'd63, 8'd14};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd164, 8'd87, 8'd43};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd140, 8'd46, 8'd20};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd160, 8'd68, 8'd27};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd154, 8'd61, 8'd18};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd151, 8'd56, 8'd12};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd162, 8'd65, 8'd22};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd182, 8'd85, 8'd43};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd188, 8'd94, 8'd58};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd163, 8'd74, 8'd42};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd130, 8'd43, 8'd13};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd177, 8'd78, 8'd39};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd184, 8'd81, 8'd40};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd180, 8'd73, 8'd29};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd173, 8'd62, 8'd17};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd189, 8'd76, 8'd32};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd186, 8'd75, 8'd32};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd165, 8'd56, 8'd17};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd176, 8'd68, 8'd32};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd193, 8'd69, 8'd35};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd162, 8'd54, 8'd18};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd153, 8'd58, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd127, 8'd33, 8'd5};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd162, 8'd56, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd195, 8'd82, 8'd52};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd184, 8'd72, 8'd32};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd170, 8'd64, 8'd16};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd156, 8'd51, 8'd6};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd183, 8'd76, 8'd34};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd179, 8'd70, 8'd29};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd169, 8'd57, 8'd19};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd188, 8'd78, 8'd41};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd195, 8'd89, 8'd50};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd184, 8'd82, 8'd44};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd148, 8'd49, 8'd10};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd139, 8'd42, 8'd7};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd178, 8'd87, 8'd56};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd158, 8'd74, 8'd48};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd117, 8'd39, 8'd17};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd91, 8'd13, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd111, 8'd27, 8'd3};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd159, 8'd68, 8'd39};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd22};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd141, 8'd41, 8'd5};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd143, 8'd50, 8'd17};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd127, 8'd41, 8'd8};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd150, 8'd61, 8'd21};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd11};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd148, 8'd52, 8'd10};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd123, 8'd37, 8'd10};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd95, 8'd22, 8'd7};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd112, 8'd37, 8'd14};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd138, 8'd54, 8'd20};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd13};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd154, 8'd59, 8'd15};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd137, 8'd49, 8'd11};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd123, 8'd41, 8'd4};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd139, 8'd54, 8'd13};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd148, 8'd56, 8'd9};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd121, 8'd43, 8'd7};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd125, 8'd77, 8'd55};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd173, 8'd163, 8'd162};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd166, 8'd185, 8'd192};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd137, 8'd161, 8'd171};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd142, 8'd165, 8'd173};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd149, 8'd167, 8'd179};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd164, 8'd183, 8'd198};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd183, 8'd161, 8'd147};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd119, 8'd88, 8'd68};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd122, 8'd76, 8'd50};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd118, 8'd56, 8'd19};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd128, 8'd51, 8'd7};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd141, 8'd53, 8'd5};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd150, 8'd54, 8'd4};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd158, 8'd58, 8'd8};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd165, 8'd69, 8'd9};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd177, 8'd81, 8'd20};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd178, 8'd83, 8'd19};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd170, 8'd70, 8'd8};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd173, 8'd63, 8'd10};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd191, 8'd71, 8'd34};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd209, 8'd79, 8'd57};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd216, 8'd78, 8'd67};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd181, 8'd39, 8'd37};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd172, 8'd28, 8'd27};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd159, 8'd13, 8'd13};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd154, 8'd4, 8'd5};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd153, 8'd3, 8'd4};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd152, 8'd6, 8'd6};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd152, 8'd8, 8'd7};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd149, 8'd10, 8'd7};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd143, 8'd0, 8'd5};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd157, 8'd4, 8'd0};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd162, 8'd16, 8'd1};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd169, 8'd30, 8'd23};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd188, 8'd28, 8'd38};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd205, 8'd26, 8'd29};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd225, 8'd83, 8'd35};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd250, 8'd168, 8'd66};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd248, 8'd166, 8'd18};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd235, 8'd149, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd182, 8'd91, 8'd8};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd142, 8'd52, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd149, 8'd68, 8'd5};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd161, 8'd91, 8'd19};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd168, 8'd109, 8'd31};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd186, 8'd133, 8'd53};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd207, 8'd154, 8'd38};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd228, 8'd179, 8'd61};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd243, 8'd201, 8'd81};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd243, 8'd209, 8'd86};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd239, 8'd209, 8'd87};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd241, 8'd211, 8'd89};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd90};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd240, 8'd210, 8'd88};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd244, 8'd206, 8'd123};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd245, 8'd209, 8'd125};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd212, 8'd130};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd250, 8'd217, 8'd138};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd252, 8'd223, 8'd145};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd152};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd157};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd160};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd183};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd185};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd188};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd191};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd194};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd197};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd200};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd202};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd212};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd213};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd212};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd202};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd190};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd250, 8'd227, 8'd177};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd169};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd247, 8'd228, 8'd169};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd233, 8'd224, 8'd167};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd236, 8'd232, 8'd185};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd91: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd242, 8'd239, 8'd186};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd233, 8'd223, 8'd136};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd227, 8'd208, 8'd105};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd232, 8'd203, 8'd101};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd244, 8'd207, 8'd118};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd134};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd238, 8'd211, 8'd108};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd240, 8'd212, 8'd112};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd240, 8'd215, 8'd115};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd241, 8'd217, 8'd119};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd241, 8'd219, 8'd120};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd240, 8'd218, 8'd119};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd239, 8'd215, 8'd117};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd238, 8'd214, 8'd116};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd249, 8'd210, 8'd115};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd249, 8'd209, 8'd113};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd110};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd249, 8'd206, 8'd102};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd250, 8'd203, 8'd97};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd251, 8'd200, 8'd91};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd251, 8'd199, 8'd87};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd250, 8'd199, 8'd84};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd247, 8'd210, 8'd96};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd247, 8'd210, 8'd96};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd249, 8'd209, 8'd95};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd249, 8'd210, 8'd93};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd249, 8'd208, 8'd90};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd88};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd88};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd251, 8'd207, 8'd86};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd243, 8'd202, 8'd84};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd243, 8'd201, 8'd83};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd241, 8'd196, 8'd81};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd234, 8'd183, 8'd74};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd223, 8'd163, 8'd65};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd210, 8'd138, 8'd54};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd198, 8'd114, 8'd44};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd192, 8'd99, 8'd38};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd178, 8'd70, 8'd31};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd159, 8'd59, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd250, 8'd167, 8'd47};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd233, 8'd164, 8'd24};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd248, 8'd176, 8'd56};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd220, 8'd118, 8'd46};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd192, 8'd41, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd225, 8'd37, 8'd51};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd179, 8'd17, 8'd15};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd169, 8'd14, 8'd12};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd157, 8'd9, 8'd5};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd144, 8'd5, 8'd0};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd137, 8'd4, 8'd0};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd137, 8'd4, 8'd0};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd139, 8'd5, 8'd2};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd142, 8'd7, 8'd4};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd155, 8'd4, 8'd11};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd172, 8'd21, 8'd26};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd196, 8'd47, 8'd49};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd212, 8'd69, 8'd65};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd213, 8'd80, 8'd65};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd200, 8'd79, 8'd48};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd181, 8'd73, 8'd27};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd168, 8'd67, 8'd13};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd179, 8'd87, 8'd10};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd184, 8'd92, 8'd15};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd185, 8'd93, 8'd18};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd175, 8'd84, 8'd13};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd158, 8'd69, 8'd3};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd146, 8'd57, 8'd1};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd140, 8'd54, 8'd5};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd140, 8'd56, 8'd12};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd110, 8'd50, 8'd16};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd129, 8'd67, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd136, 8'd82, 8'd46};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd128, 8'd96, 8'd73};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd156, 8'd153, 8'd146};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd161, 8'd179, 8'd183};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd166, 8'd186, 8'd193};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd162, 8'd181, 8'd185};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd146, 8'd150, 8'd161};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd136, 8'd155, 8'd159};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd146, 8'd147, 8'd142};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd144, 8'd88, 8'd75};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd140, 8'd53, 8'd23};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd137, 8'd56, 8'd9};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd165, 8'd86, 8'd43};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd150, 8'd55, 8'd25};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd163, 8'd67, 8'd25};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd13};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd153, 8'd55, 8'd10};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd164, 8'd63, 8'd19};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd177, 8'd78, 8'd36};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd187, 8'd91, 8'd53};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd170, 8'd77, 8'd44};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd138, 8'd49, 8'd19};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd175, 8'd76, 8'd37};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd188, 8'd85, 8'd44};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd181, 8'd74, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd176, 8'd65, 8'd20};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd189, 8'd76, 8'd32};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd183, 8'd72, 8'd29};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd167, 8'd58, 8'd19};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd178, 8'd70, 8'd34};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd195, 8'd68, 8'd33};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd170, 8'd60, 8'd25};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd156, 8'd59, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd128, 8'd33, 8'd3};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd164, 8'd59, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd194, 8'd79, 8'd48};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd187, 8'd74, 8'd34};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd176, 8'd68, 8'd21};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd167, 8'd60, 8'd16};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd172, 8'd63, 8'd20};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd181, 8'd69, 8'd29};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd171, 8'd58, 8'd18};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd184, 8'd72, 8'd34};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd175, 8'd67, 8'd29};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd183, 8'd79, 8'd40};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd174, 8'd75, 8'd34};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd129, 8'd38, 8'd11};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd124, 8'd40, 8'd16};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd162, 8'd89, 8'd70};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd119, 8'd53, 8'd37};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd61, 8'd0, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd112, 8'd36, 8'd12};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd160, 8'd71, 8'd39};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd158, 8'd60, 8'd23};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd141, 8'd41, 8'd7};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd142, 8'd49, 8'd16};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd126, 8'd40, 8'd7};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd149, 8'd59, 8'd22};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd13};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd147, 8'd51, 8'd11};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd122, 8'd36, 8'd9};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd95, 8'd22, 8'd7};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd110, 8'd38, 8'd16};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd140, 8'd55, 8'd24};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd13};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd13};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd137, 8'd49, 8'd11};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd128, 8'd44, 8'd7};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd144, 8'd55, 8'd13};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd148, 8'd52, 8'd4};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd117, 8'd39, 8'd3};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd126, 8'd79, 8'd59};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd172, 8'd164, 8'd162};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd160, 8'd178, 8'd188};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd132, 8'd159, 8'd170};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd141, 8'd163, 8'd174};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd143, 8'd162, 8'd176};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd159, 8'd178, 8'd195};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd181, 8'd159, 8'd148};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd115, 8'd82, 8'd65};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd117, 8'd70, 8'd42};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd116, 8'd51, 8'd13};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd131, 8'd50, 8'd3};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd145, 8'd55, 8'd3};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd148, 8'd54, 8'd2};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd4};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd174, 8'd73, 8'd17};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd169, 8'd68, 8'd12};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd166, 8'd61, 8'd6};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd174, 8'd62, 8'd14};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd195, 8'd75, 8'd40};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd214, 8'd84, 8'd62};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd210, 8'd71, 8'd64};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd197, 8'd53, 8'd53};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd162, 8'd20, 8'd19};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd155, 8'd13, 8'd12};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd147, 8'd3, 8'd3};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd142, 8'd0, 8'd0};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd142, 8'd0, 8'd0};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd146, 8'd1, 8'd0};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd152, 8'd7, 8'd4};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd155, 8'd10, 8'd7};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd151, 8'd0, 8'd7};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd168, 8'd9, 8'd5};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd177, 8'd23, 8'd11};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd185, 8'd38, 8'd31};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd199, 8'd33, 8'd43};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd209, 8'd29, 8'd32};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd226, 8'd86, 8'd37};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd250, 8'd171, 8'd66};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd247, 8'd165, 8'd21};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd240, 8'd151, 8'd35};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd193, 8'd97, 8'd20};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd154, 8'd58, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd160, 8'd72, 8'd9};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd168, 8'd94, 8'd21};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd174, 8'd113, 8'd32};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd191, 8'd139, 8'd55};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd226, 8'd164, 8'd65};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd245, 8'd188, 8'd85};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd102};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd101};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd252, 8'd211, 8'd93};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd252, 8'd212, 8'd90};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd252, 8'd211, 8'd87};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd252, 8'd208, 8'd83};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd249, 8'd207, 8'd71};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd72};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd248, 8'd208, 8'd74};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd247, 8'd209, 8'd76};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd246, 8'd209, 8'd77};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd247, 8'd210, 8'd80};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd245, 8'd210, 8'd80};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd245, 8'd210, 8'd82};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd251, 8'd209, 8'd89};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd90};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd249, 8'd208, 8'd92};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd248, 8'd208, 8'd95};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd246, 8'd208, 8'd99};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd245, 8'd208, 8'd101};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd242, 8'd208, 8'd101};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd242, 8'd207, 8'd103};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd227, 8'd214, 8'd86};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd227, 8'd207, 8'd92};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd230, 8'd205, 8'd104};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd241, 8'd207, 8'd117};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd248, 8'd213, 8'd119};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd245, 8'd215, 8'd105};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd231, 8'd207, 8'd75};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd219, 8'd198, 8'd53};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd237, 8'd227, 8'd155};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd241, 8'd234, 8'd179};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd92: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd254, 8'd241, 8'd189};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd234, 8'd213, 8'd134};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd228, 8'd196, 8'd93};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd202, 8'd78};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd80};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd252, 8'd214, 8'd79};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd250, 8'd212, 8'd77};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd247, 8'd209, 8'd74};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd244, 8'd206, 8'd73};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd240, 8'd203, 8'd71};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd235, 8'd202, 8'd71};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd232, 8'd202, 8'd72};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd231, 8'd202, 8'd74};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd245, 8'd201, 8'd76};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd247, 8'd202, 8'd75};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd251, 8'd203, 8'd75};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd254, 8'd205, 8'd74};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd73};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd74};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd72};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd73};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd253, 8'd212, 8'd84};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd253, 8'd212, 8'd84};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd84};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd86};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd86};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd88};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd90};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd90};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd253, 8'd215, 8'd108};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd106};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd243, 8'd201, 8'd99};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd230, 8'd184, 8'd90};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd214, 8'd156, 8'd74};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd195, 8'd124, 8'd58};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd178, 8'd97, 8'd44};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd168, 8'd79, 8'd35};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd188, 8'd76, 8'd36};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd168, 8'd68, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd53};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd237, 8'd177, 8'd31};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd249, 8'd185, 8'd59};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd221, 8'd121, 8'd45};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd194, 8'd42, 8'd21};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd230, 8'd38, 8'd51};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd193, 8'd27, 8'd27};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd185, 8'd23, 8'd21};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd169, 8'd16, 8'd11};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd156, 8'd8, 8'd4};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd145, 8'd3, 8'd0};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd140, 8'd3, 8'd0};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd138, 8'd3, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd139, 8'd4, 8'd0};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd156, 8'd5, 8'd10};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd155, 8'd4, 8'd11};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd165, 8'd14, 8'd21};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd191, 8'd42, 8'd44};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd216, 8'd74, 8'd70};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd222, 8'd90, 8'd75};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd206, 8'd85, 8'd58};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd186, 8'd72, 8'd38};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd176, 8'd76, 8'd14};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd181, 8'd83, 8'd20};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd184, 8'd91, 8'd24};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd178, 8'd89, 8'd23};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd163, 8'd78, 8'd14};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd149, 8'd64, 8'd7};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd141, 8'd55, 8'd4};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd138, 8'd52, 8'd5};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd117, 8'd55, 8'd16};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd121, 8'd58, 8'd17};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd132, 8'd74, 8'd36};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd136, 8'd99, 8'd73};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd166, 8'd157, 8'd150};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd166, 8'd179, 8'd185};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd159, 8'd182, 8'd188};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd149, 8'd170, 8'd173};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd184, 8'd191, 8'd199};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd170, 8'd191, 8'd192};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd159, 8'd160, 8'd155};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd149, 8'd92, 8'd83};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd130, 8'd43, 8'd16};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd131, 8'd49, 8'd2};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd170, 8'd89, 8'd44};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd162, 8'd63, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd164, 8'd65, 8'd23};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd154, 8'd53, 8'd9};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd158, 8'd55, 8'd10};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd170, 8'd65, 8'd20};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd177, 8'd74, 8'd33};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd87, 8'd48};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd175, 8'd78, 8'd45};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd142, 8'd47, 8'd17};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd174, 8'd75, 8'd36};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd191, 8'd88, 8'd47};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd182, 8'd75, 8'd31};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd179, 8'd68, 8'd23};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd190, 8'd77, 8'd33};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd180, 8'd69, 8'd26};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd170, 8'd61, 8'd22};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd180, 8'd72, 8'd36};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd194, 8'd67, 8'd32};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd180, 8'd68, 8'd31};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd157, 8'd60, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd131, 8'd34, 8'd2};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd168, 8'd60, 8'd32};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd193, 8'd76, 8'd43};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd191, 8'd75, 8'd34};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd182, 8'd74, 8'd25};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd175, 8'd68, 8'd22};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd164, 8'd56, 8'd10};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd179, 8'd66, 8'd24};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd175, 8'd62, 8'd22};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd185, 8'd72, 8'd32};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd172, 8'd63, 8'd24};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd178, 8'd75, 8'd34};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd181, 8'd79, 8'd39};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd176, 8'd82, 8'd57};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd102, 8'd20, 8'd0};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd109, 8'd42, 8'd26};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd106, 8'd50, 8'd37};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd80, 8'd23, 8'd6};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd108, 8'd38, 8'd13};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd143, 8'd57, 8'd24};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd165, 8'd66, 8'd27};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd140, 8'd40, 8'd6};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd142, 8'd49, 8'd18};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd126, 8'd39, 8'd9};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd149, 8'd59, 8'd22};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd13};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd147, 8'd51, 8'd11};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd122, 8'd36, 8'd11};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd94, 8'd20, 8'd7};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd111, 8'd38, 8'd19};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd141, 8'd58, 8'd28};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd15};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd150, 8'd53, 8'd10};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd138, 8'd49, 8'd9};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd133, 8'd48, 8'd11};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd149, 8'd58, 8'd14};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd148, 8'd48, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd118, 8'd42, 8'd8};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd137, 8'd90, 8'd72};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd177, 8'd171, 8'd171};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd160, 8'd180, 8'd191};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd135, 8'd163, 8'd174};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd145, 8'd169, 8'd179};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd144, 8'd166, 8'd179};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd160, 8'd181, 8'd200};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd179, 8'd155, 8'd143};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd110, 8'd75, 8'd56};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd116, 8'd65, 8'd34};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd123, 8'd54, 8'd12};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd138, 8'd55, 8'd5};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd143, 8'd53, 8'd1};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd149, 8'd57, 8'd8};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd176, 8'd74, 8'd25};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd165, 8'd58, 8'd12};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd169, 8'd56, 8'd16};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd198, 8'd75, 8'd44};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd223, 8'd92, 8'd72};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd222, 8'd83, 8'd76};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd197, 8'd52, 8'd55};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd173, 8'd27, 8'd37};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd154, 8'd11, 8'd13};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd150, 8'd7, 8'd9};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd143, 8'd1, 8'd0};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd137, 8'd0, 8'd0};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd137, 8'd0, 8'd0};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd145, 8'd0, 8'd0};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd154, 8'd5, 8'd1};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd162, 8'd10, 8'd7};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd167, 8'd10, 8'd17};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd187, 8'd19, 8'd18};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd197, 8'd35, 8'd24};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd201, 8'd46, 8'd41};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd209, 8'd38, 8'd47};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd215, 8'd31, 8'd33};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd229, 8'd89, 8'd38};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd252, 8'd178, 8'd71};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd245, 8'd168, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd50};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd203, 8'd104, 8'd36};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd160, 8'd58, 8'd10};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd156, 8'd60, 8'd10};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd158, 8'd77, 8'd14};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd166, 8'd98, 8'd27};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd187, 8'd129, 8'd56};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd212, 8'd154, 8'd70};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd233, 8'd179, 8'd91};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd252, 8'd203, 8'd111};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd254, 8'd212, 8'd112};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd252, 8'd213, 8'd108};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd109};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd107};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd104};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd98};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd97};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd95};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd252, 8'd216, 8'd94};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd249, 8'd213, 8'd91};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd246, 8'd211, 8'd91};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd244, 8'd209, 8'd89};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd243, 8'd208, 8'd88};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd249, 8'd210, 8'd71};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd248, 8'd210, 8'd73};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd76};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd78};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd249, 8'd212, 8'd80};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd249, 8'd212, 8'd82};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd248, 8'd213, 8'd85};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd248, 8'd213, 8'd85};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd236, 8'd205, 8'd65};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd248, 8'd216, 8'd73};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd78};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd73};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd245, 8'd210, 8'd66};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd236, 8'd204, 8'd67};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd238, 8'd211, 8'd80};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd244, 8'd220, 8'd94};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd187};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd254, 8'd245, 8'd204};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd93: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd206};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd253, 8'd227, 8'd153};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd242, 8'd210, 8'd99};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd235, 8'd199, 8'd63};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd247, 8'd215, 8'd92};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd253, 8'd219, 8'd95};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd102};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd107};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd108};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd110};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd246, 8'd223, 8'd107};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd239, 8'd219, 8'd106};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd243, 8'd217, 8'd106};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd241, 8'd218, 8'd106};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd241, 8'd218, 8'd106};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd241, 8'd218, 8'd104};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd240, 8'd217, 8'd103};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd240, 8'd217, 8'd101};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd240, 8'd217, 8'd101};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd239, 8'd217, 8'd98};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd251, 8'd220, 8'd103};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd103};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd103};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd253, 8'd218, 8'd102};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd253, 8'd218, 8'd102};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd253, 8'd216, 8'd101};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd101};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd101};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd254, 8'd224, 8'd114};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd110};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd242, 8'd208, 8'd101};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd231, 8'd189, 8'd87};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd214, 8'd160, 8'd70};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd195, 8'd128, 8'd50};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd177, 8'd98, 8'd32};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd167, 8'd81, 8'd24};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd188, 8'd73, 8'd29};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd171, 8'd70, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd188, 8'd60};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd244, 8'd190, 8'd38};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd253, 8'd196, 8'd65};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd224, 8'd129, 8'd49};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd199, 8'd47, 8'd23};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd238, 8'd42, 8'd52};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd209, 8'd41, 8'd40};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd200, 8'd35, 8'd33};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd187, 8'd25, 8'd23};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd170, 8'd15, 8'd11};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd157, 8'd8, 8'd4};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd149, 8'd4, 8'd1};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd145, 8'd3, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd145, 8'd3, 8'd1};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd160, 8'd7, 8'd10};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd154, 8'd1, 8'd4};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd154, 8'd0, 8'd5};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd169, 8'd15, 8'd23};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd193, 8'd44, 8'd46};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd215, 8'd73, 8'd69};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd222, 8'd90, 8'd77};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd222, 8'd95, 8'd76};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd179, 8'd72, 8'd26};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd180, 8'd78, 8'd29};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd182, 8'd87, 8'd31};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd180, 8'd91, 8'd33};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd172, 8'd88, 8'd28};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd157, 8'd75, 8'd19};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd141, 8'd58, 8'd8};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd132, 8'd46, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd125, 8'd58, 8'd15};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd121, 8'd53, 8'd6};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd130, 8'd65, 8'd23};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd138, 8'd93, 8'd64};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd168, 8'd151, 8'd141};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd171, 8'd181, 8'd183};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd169, 8'd190, 8'd193};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd154, 8'd175, 8'd176};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd211, 8'd220, 8'd225};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd183, 8'd207, 8'd207};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd147, 8'd149, 8'd146};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd138, 8'd83, 8'd76};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd126, 8'd36, 8'd12};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd133, 8'd49, 8'd5};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd169, 8'd86, 8'd42};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd154, 8'd54, 8'd20};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd166, 8'd63, 8'd22};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd156, 8'd50, 8'd8};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd165, 8'd58, 8'd14};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd177, 8'd68, 8'd25};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd178, 8'd71, 8'd29};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd82, 8'd45};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd175, 8'd75, 8'd43};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd139, 8'd41, 8'd12};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd172, 8'd73, 8'd34};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd194, 8'd91, 8'd50};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd183, 8'd76, 8'd32};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd182, 8'd71, 8'd26};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd190, 8'd77, 8'd33};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd177, 8'd66, 8'd23};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd172, 8'd63, 8'd24};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd182, 8'd74, 8'd38};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd195, 8'd67, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd187, 8'd75, 8'd37};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd159, 8'd61, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd131, 8'd34, 8'd2};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd171, 8'd62, 8'd33};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd191, 8'd74, 8'd41};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd193, 8'd78, 8'd34};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd190, 8'd80, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd176, 8'd68, 8'd22};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd165, 8'd54, 8'd9};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd178, 8'd65, 8'd21};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd177, 8'd61, 8'd20};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd185, 8'd72, 8'd32};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd190, 8'd81, 8'd40};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd180, 8'd74, 8'd34};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd160, 8'd59, 8'd17};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd194, 8'd92, 8'd67};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd159, 8'd71, 8'd49};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd82, 8'd16, 8'd0};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd74, 8'd22, 8'd9};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd94, 8'd42, 8'd28};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd100, 8'd36, 8'd11};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd138, 8'd54, 8'd20};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd162, 8'd63, 8'd22};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd140, 8'd40, 8'd8};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd125, 8'd38, 8'd10};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd148, 8'd58, 8'd23};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd13};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd146, 8'd50, 8'd12};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd121, 8'd35, 8'd12};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd94, 8'd20, 8'd9};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd110, 8'd39, 8'd21};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd142, 8'd58, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd148, 8'd51, 8'd9};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd140, 8'd48, 8'd9};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd140, 8'd50, 8'd13};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd154, 8'd59, 8'd15};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd146, 8'd44, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd115, 8'd39, 8'd7};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd138, 8'd93, 8'd74};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd176, 8'd170, 8'd172};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd152, 8'd174, 8'd185};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd132, 8'd160, 8'd172};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd144, 8'd168, 8'd180};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd139, 8'd161, 8'd175};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd154, 8'd177, 8'd195};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd170, 8'd147, 8'd131};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd108, 8'd72, 8'd48};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd124, 8'd70, 8'd34};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd134, 8'd61, 8'd16};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd146, 8'd60, 8'd9};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd145, 8'd53, 8'd4};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd141, 8'd50, 8'd5};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd145, 8'd56, 8'd14};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd170, 8'd68, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd173, 8'd64, 8'd31};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd191, 8'd73, 8'd47};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd217, 8'd90, 8'd73};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd224, 8'd87, 8'd79};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd202, 8'd59, 8'd61};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd175, 8'd30, 8'd37};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd162, 8'd16, 8'd27};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd150, 8'd7, 8'd13};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd147, 8'd7, 8'd10};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd143, 8'd3, 8'd4};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd138, 8'd0, 8'd0};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd138, 8'd0, 8'd0};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd147, 8'd0, 8'd0};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd160, 8'd8, 8'd3};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd171, 8'd16, 8'd11};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd190, 8'd26, 8'd35};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd208, 8'd34, 8'd33};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd217, 8'd46, 8'd36};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd216, 8'd52, 8'd50};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd217, 8'd39, 8'd51};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd218, 8'd32, 8'd33};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd231, 8'd94, 8'd40};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd75};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd243, 8'd174, 8'd35};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd245, 8'd164, 8'd57};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd207, 8'd109, 8'd44};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd166, 8'd59, 8'd17};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd160, 8'd57, 8'd16};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd165, 8'd73, 8'd22};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd178, 8'd99, 8'd42};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd204, 8'd134, 8'd75};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd212, 8'd157, 8'd67};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd232, 8'd181, 8'd89};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd249, 8'd207, 8'd109};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd249, 8'd214, 8'd112};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd247, 8'd216, 8'd110};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd248, 8'd220, 8'd111};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd250, 8'd222, 8'd112};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd108};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd250, 8'd225, 8'd107};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd250, 8'd225, 8'd107};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd249, 8'd224, 8'd106};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd248, 8'd223, 8'd105};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd247, 8'd222, 8'd104};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd246, 8'd221, 8'd103};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd102};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd246, 8'd219, 8'd102};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd240, 8'd224, 8'd111};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd240, 8'd224, 8'd111};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd242, 8'd224, 8'd112};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd245, 8'd225, 8'd113};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd247, 8'd225, 8'd114};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd249, 8'd227, 8'd116};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd251, 8'd227, 8'd117};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd251, 8'd227, 8'd117};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd136};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd119};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd86};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd250, 8'd212, 8'd51};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd222, 8'd192, 8'd42};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd220, 8'd194, 8'd84};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd245, 8'd220, 8'd163};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd94: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd219};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd247, 8'd222, 8'd166};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd228, 8'd200, 8'd127};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd218, 8'd170, 8'd68};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd225, 8'd176, 8'd73};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd238, 8'd187, 8'd80};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd251, 8'd198, 8'd92};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd105};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd117};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd127};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd254, 8'd223, 8'd133};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd150};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd151};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd150};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd254, 8'd236, 8'd150};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd251, 8'd236, 8'd151};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd247, 8'd237, 8'd152};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd244, 8'd236, 8'd153};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd244, 8'd236, 8'd153};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd146};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd254, 8'd237, 8'd145};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd144};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd253, 8'd233, 8'd144};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd252, 8'd231, 8'd142};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd252, 8'd228, 8'd140};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd250, 8'd226, 8'd140};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd250, 8'd226, 8'd140};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd251, 8'd223, 8'd124};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd249, 8'd220, 8'd120};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd245, 8'd210, 8'd110};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd235, 8'd191, 8'd92};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd221, 8'd164, 8'd74};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd205, 8'd133, 8'd51};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd192, 8'd104, 8'd33};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd182, 8'd87, 8'd23};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd179, 8'd60, 8'd17};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd166, 8'd65, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd61};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd247, 8'd201, 8'd45};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd73};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd232, 8'd140, 8'd57};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd210, 8'd56, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd251, 8'd51, 8'd61};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd54, 8'd53};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd214, 8'd46, 8'd45};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd199, 8'd34, 8'd32};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd185, 8'd21, 8'd20};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd170, 8'd10, 8'd10};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd161, 8'd6, 8'd4};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd156, 8'd4, 8'd3};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd153, 8'd3, 8'd2};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd156, 8'd4, 8'd3};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd157, 8'd3, 8'd5};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd157, 8'd2, 8'd8};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd161, 8'd4, 8'd13};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd172, 8'd19, 8'd24};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd193, 8'd44, 8'd46};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd218, 8'd76, 8'd72};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd235, 8'd98, 8'd88};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd202, 8'd89, 8'd57};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd189, 8'd83, 8'd44};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd174, 8'd77, 8'd32};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd165, 8'd77, 8'd27};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd163, 8'd80, 8'd26};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd158, 8'd77, 8'd24};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd148, 8'd64, 8'd17};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd140, 8'd53, 8'd8};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd139, 8'd69, 8'd18};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd141, 8'd65, 8'd15};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd144, 8'd72, 8'd24};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd132, 8'd79, 8'd47};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd151, 8'd129, 8'd116};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd167, 8'd171, 8'd170};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd178, 8'd196, 8'd196};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd163, 8'd183, 8'd181};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd194, 8'd205, 8'd207};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd172, 8'd198, 8'd195};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd134, 8'd139, 8'd135};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd140, 8'd85, 8'd80};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd129, 8'd38, 8'd17};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd137, 8'd53, 8'd9};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd169, 8'd85, 8'd39};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd148, 8'd45, 8'd10};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd167, 8'd61, 8'd19};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd157, 8'd50, 8'd6};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd174, 8'd63, 8'd18};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd187, 8'd74, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd182, 8'd70, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd78, 8'd40};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd173, 8'd70, 8'd37};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd133, 8'd32, 8'd2};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd171, 8'd72, 8'd33};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd197, 8'd94, 8'd53};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd183, 8'd76, 8'd32};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd184, 8'd73, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd78, 8'd34};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd174, 8'd63, 8'd20};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd174, 8'd65, 8'd26};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd183, 8'd75, 8'd39};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd195, 8'd66, 8'd27};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd193, 8'd79, 8'd42};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd159, 8'd61, 8'd24};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd132, 8'd33, 8'd1};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd172, 8'd63, 8'd34};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd190, 8'd71, 8'd37};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd196, 8'd79, 8'd36};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd195, 8'd83, 8'd33};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd178, 8'd70, 8'd23};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd171, 8'd60, 8'd14};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd182, 8'd67, 8'd23};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd179, 8'd62, 8'd19};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd175, 8'd59, 8'd18};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd198, 8'd86, 8'd46};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd179, 8'd72, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd156, 8'd53, 8'd12};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd175, 8'd62, 8'd32};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd195, 8'd101, 8'd75};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd121, 8'd53, 8'd34};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd66, 8'd17, 8'd3};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd77, 8'd31, 8'd15};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd104, 8'd44, 8'd20};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd144, 8'd61, 8'd27};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd157, 8'd60, 8'd18};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd140, 8'd40, 8'd8};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd125, 8'd38, 8'd10};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd148, 8'd58, 8'd24};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd14};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd146, 8'd49, 8'd14};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd121, 8'd35, 8'd12};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd93, 8'd19, 8'd8};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd111, 8'd39, 8'd24};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd144, 8'd60, 8'd34};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd147, 8'd48, 8'd7};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd9};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd146, 8'd54, 8'd17};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd157, 8'd60, 8'd15};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd147, 8'd41, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd112, 8'd37, 8'd5};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd141, 8'd95, 8'd79};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd176, 8'd172, 8'd173};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd149, 8'd171, 8'd184};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd130, 8'd160, 8'd171};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd142, 8'd169, 8'd180};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd136, 8'd159, 8'd173};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd151, 8'd173, 8'd194};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd158, 8'd134, 8'd110};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd113, 8'd77, 8'd45};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd139, 8'd81, 8'd41};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd143, 8'd67, 8'd17};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd150, 8'd60, 8'd8};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd12};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd143, 8'd54, 8'd14};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd140, 8'd51, 8'd17};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd171, 8'd70, 8'd42};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd188, 8'd79, 8'd56};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd209, 8'd89, 8'd75};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd214, 8'd82, 8'd77};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd199, 8'd59, 8'd60};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd175, 8'd32, 8'd38};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd159, 8'd15, 8'd24};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd152, 8'd11, 8'd19};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd147, 8'd4, 8'd10};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd146, 8'd5, 8'd11};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd145, 8'd7, 8'd7};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd141, 8'd3, 8'd1};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd141, 8'd2, 8'd0};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd154, 8'd6, 8'd2};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd172, 8'd19, 8'd13};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd188, 8'd29, 8'd25};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd210, 8'd43, 8'd51};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd229, 8'd49, 8'd50};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd234, 8'd57, 8'd49};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd226, 8'd58, 8'd55};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd222, 8'd40, 8'd52};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd221, 8'd33, 8'd34};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd234, 8'd97, 8'd43};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd81};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd247, 8'd190, 8'd38};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd244, 8'd172, 8'd52};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd202, 8'd108, 8'd34};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd163, 8'd55, 8'd8};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd165, 8'd56, 8'd13};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd177, 8'd75, 8'd27};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd189, 8'd99, 8'd46};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd211, 8'd132, 8'd76};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd232, 8'd170, 8'd83};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd250, 8'd195, 8'd105};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd128};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd132};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd132};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd136};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd137};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd254, 8'd227, 8'd136};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd253, 8'd234, 8'd132};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd253, 8'd234, 8'd132};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd131};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd131};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd131};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd129};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd129};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd129};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd154};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd150};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd146};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd140};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd132};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd125};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd120};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd254, 8'd211, 8'd119};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd105};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd238, 8'd173, 8'd73};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd214, 8'd157, 8'd44};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd210, 8'd167, 8'd54};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd229, 8'd198, 8'd108};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd248, 8'd228, 8'd178};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd95: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd89};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd253, 8'd173, 8'd76};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd239, 8'd157, 8'd57};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd230, 8'd146, 8'd47};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd228, 8'd148, 8'd49};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd235, 8'd162, 8'd68};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd246, 8'd180, 8'd94};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd254, 8'd193, 8'd112};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd251, 8'd208, 8'd129};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd252, 8'd211, 8'd132};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd217, 8'd139};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd149};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd159};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd170};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd176};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd180};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd249, 8'd242, 8'd170};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd249, 8'd242, 8'd170};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd249, 8'd241, 8'd169};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd248, 8'd239, 8'd170};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd249, 8'd239, 8'd170};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd250, 8'd236, 8'd171};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd249, 8'd235, 8'd170};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd249, 8'd235, 8'd170};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd147};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd219, 8'd141};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd249, 8'd206, 8'd127};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd237, 8'd184, 8'd104};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd221, 8'd153, 8'd78};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd203, 8'd118, 8'd51};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd188, 8'd88, 8'd29};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd179, 8'd69, 8'd16};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd171, 8'd50, 8'd7};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd160, 8'd60, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd59};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd206, 8'd49};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd79};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd238, 8'd147, 8'd64};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd218, 8'd64, 8'd38};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd59, 8'd69};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd230, 8'd62, 8'd59};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd222, 8'd54, 8'd53};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd209, 8'd39, 8'd39};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd193, 8'd25, 8'd25};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd179, 8'd13, 8'd13};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd169, 8'd6, 8'd7};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd162, 8'd4, 8'd5};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd159, 8'd3, 8'd4};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd150, 8'd0, 8'd0};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd157, 8'd3, 8'd3};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd163, 8'd7, 8'd11};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd164, 8'd7, 8'd14};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd167, 8'd12, 8'd20};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd180, 8'd30, 8'd32};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd204, 8'd58, 8'd58};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd223, 8'd81, 8'd77};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd228, 8'd112, 8'd87};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd200, 8'd91, 8'd62};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd165, 8'd67, 8'd28};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd147, 8'd59, 8'd13};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd148, 8'd66, 8'd16};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd156, 8'd74, 8'd24};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd157, 8'd73, 8'd27};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd156, 8'd69, 8'd26};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd156, 8'd83, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd165, 8'd86, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd161, 8'd85, 8'd35};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd127, 8'd68, 8'd34};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd133, 8'd105, 8'd91};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd159, 8'd159, 8'd157};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd181, 8'd197, 8'd196};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd164, 8'd183, 8'd177};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd187, 8'd201, 8'd201};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd175, 8'd204, 8'd200};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd144, 8'd148, 8'd147};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd152, 8'd97, 8'd94};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd133, 8'd42, 8'd21};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd137, 8'd52, 8'd11};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd174, 8'd87, 8'd42};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd157, 8'd54, 8'd19};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd167, 8'd60, 8'd18};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd158, 8'd49, 8'd6};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd178, 8'd65, 8'd21};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd191, 8'd78, 8'd34};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd183, 8'd70, 8'd28};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd185, 8'd75, 8'd38};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd171, 8'd66, 8'd34};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd130, 8'd26, 8'd0};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd170, 8'd71, 8'd32};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd198, 8'd95, 8'd54};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd184, 8'd77, 8'd33};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd185, 8'd74, 8'd29};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd78, 8'd34};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd173, 8'd62, 8'd19};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd175, 8'd66, 8'd27};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd184, 8'd76, 8'd40};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd195, 8'd66, 8'd27};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd196, 8'd82, 8'd45};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd161, 8'd61, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd133, 8'd34, 8'd2};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd173, 8'd64, 8'd33};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd189, 8'd70, 8'd36};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd196, 8'd79, 8'd36};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd197, 8'd85, 8'd35};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd185, 8'd74, 8'd28};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd177, 8'd65, 8'd19};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd185, 8'd70, 8'd26};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd182, 8'd65, 8'd22};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd159, 8'd43, 8'd2};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd185, 8'd73, 8'd33};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd175, 8'd68, 8'd26};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd172, 8'd69, 8'd26};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd167, 8'd47, 8'd13};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd169, 8'd70, 8'd41};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd158, 8'd87, 8'd67};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd88, 8'd41, 8'd25};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd67, 8'd24, 8'd7};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd117, 8'd59, 8'd35};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd142, 8'd62, 8'd29};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd159, 8'd61, 8'd22};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd139, 8'd38, 8'd8};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd125, 8'd38, 8'd10};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd148, 8'd58, 8'd24};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd14};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd146, 8'd49, 8'd14};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd121, 8'd35, 8'd12};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd93, 8'd19, 8'd8};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd109, 8'd40, 8'd25};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd144, 8'd60, 8'd34};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd151, 8'd55, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd146, 8'd47, 8'd6};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd9};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd147, 8'd55, 8'd16};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd159, 8'd61, 8'd16};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd146, 8'd40, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd121, 8'd46, 8'd14};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd151, 8'd108, 8'd91};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd187, 8'd183, 8'd184};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd158, 8'd180, 8'd193};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd140, 8'd169, 8'd183};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd152, 8'd178, 8'd191};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd145, 8'd168, 8'd184};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd160, 8'd182, 8'd203};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd147, 8'd123, 8'd95};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd118, 8'd82, 8'd46};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd150, 8'd93, 8'd48};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd146, 8'd69, 8'd17};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd148, 8'd58, 8'd6};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd156, 8'd63, 8'd19};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd147, 8'd57, 8'd22};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd134, 8'd47, 8'd19};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd179, 8'd79, 8'd56};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd199, 8'd92, 8'd76};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd213, 8'd92, 8'd84};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd198, 8'd65, 8'd66};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd176, 8'd35, 8'd41};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd162, 8'd18, 8'd27};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd151, 8'd10, 8'd16};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd144, 8'd5, 8'd10};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd144, 8'd0, 8'd9};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd145, 8'd4, 8'd10};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd144, 8'd8, 8'd10};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd142, 8'd7, 8'd4};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd146, 8'd7, 8'd2};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd161, 8'd14, 8'd7};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd182, 8'd27, 8'd22};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd200, 8'd38, 8'd33};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd223, 8'd53, 8'd62};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd241, 8'd59, 8'd58};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd242, 8'd63, 8'd56};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd233, 8'd61, 8'd59};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd225, 8'd41, 8'd53};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd221, 8'd33, 8'd34};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd235, 8'd100, 8'd45};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd84};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd41};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd48};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd194, 8'd104, 8'd18};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd151, 8'd44, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd156, 8'd44, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd166, 8'd60, 8'd8};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd172, 8'd77, 8'd21};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd187, 8'd102, 8'd47};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd215, 8'd142, 8'd73};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd235, 8'd168, 8'd98};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd252, 8'd195, 8'd124};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd253, 8'd206, 8'd136};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd250, 8'd211, 8'd144};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd252, 8'd218, 8'd154};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd161};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd161};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd182};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd181};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd180};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd179};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd175};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd172};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd171};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd171};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd133};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd127};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd251, 8'd194, 8'd117};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd244, 8'd181, 8'd101};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd236, 8'd168, 8'd83};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd230, 8'd156, 8'd69};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd225, 8'd145, 8'd56};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd222, 8'd141, 8'd50};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd220, 8'd150, 8'd2};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd228, 8'd160, 8'd33};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd243, 8'd179, 8'd89};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd153};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd207};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd96: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd245, 8'd230, 8'd211};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd231, 8'd206, 8'd142};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd225, 8'd183, 8'd73};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd231, 8'd165, 8'd25};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd244, 8'd150, 8'd0};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd139, 8'd0};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd130, 8'd0};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd255, 8'd131, 8'd26};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd253, 8'd128, 8'd20};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd245, 8'd125, 8'd15};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd236, 8'd121, 8'd12};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd231, 8'd122, 8'd17};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd231, 8'd124, 8'd28};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd233, 8'd129, 8'd42};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd234, 8'd131, 8'd52};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd247, 8'd141, 8'd41};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd250, 8'd141, 8'd46};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd141, 8'd53};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd57};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd254, 8'd139, 8'd56};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd248, 8'd136, 8'd50};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd239, 8'd135, 8'd40};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd235, 8'd133, 8'd33};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd238, 8'd122, 8'd39};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd234, 8'd119, 8'd38};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd226, 8'd115, 8'd36};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd217, 8'd105, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd91, 8'd24};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd201, 8'd75, 8'd16};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd196, 8'd60, 8'd8};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd194, 8'd52, 8'd4};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd191, 8'd34, 8'd3};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd193, 8'd75, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd45};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd238, 8'd224, 8'd40};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd234, 8'd221, 8'd67};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd236, 8'd169, 8'd80};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd222, 8'd73, 8'd43};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd63, 8'd66};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd245, 8'd67, 8'd67};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd248, 8'd70, 8'd70};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd244, 8'd68, 8'd68};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd232, 8'd56, 8'd56};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd211, 8'd37, 8'd36};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd193, 8'd19, 8'd18};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd182, 8'd10, 8'd8};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd179, 8'd7, 8'd5};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd169, 8'd1, 8'd0};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd163, 8'd0, 8'd0};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd158, 8'd0, 8'd0};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd158, 8'd0, 8'd0};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd164, 8'd5, 8'd1};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd177, 8'd20, 8'd15};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd190, 8'd35, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd200, 8'd45, 8'd40};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd231, 8'd80, 8'd89};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd242, 8'd111, 8'd103};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd186, 8'd77, 8'd54};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd152, 8'd52, 8'd26};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd157, 8'd55, 8'd33};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd149, 8'd45, 8'd18};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd145, 8'd49, 8'd1};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd138, 8'd53, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd139, 8'd57, 8'd9};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd158, 8'd63, 8'd35};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd174, 8'd75, 8'd43};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd155, 8'd76, 8'd17};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd117, 8'd71, 8'd19};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd146, 8'd128, 8'd118};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd178, 8'd177, 8'd193};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd180, 8'd190, 8'd200};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd200, 8'd202, 8'd214};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd186, 8'd197, 8'd203};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd150, 8'd159, 8'd154};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd132, 8'd110, 8'd89};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd118, 8'd52, 8'd17};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd133, 8'd38, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd172, 8'd77, 8'd33};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd145, 8'd62, 8'd20};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd156, 8'd56, 8'd6};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd150, 8'd53, 8'd8};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd164, 8'd67, 8'd25};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd181, 8'd75, 8'd33};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd189, 8'd77, 8'd31};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd199, 8'd87, 8'd47};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd168, 8'd70, 8'd45};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd104, 8'd21, 8'd7};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd154, 8'd69, 8'd48};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd185, 8'd87, 8'd52};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd175, 8'd60, 8'd15};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd200, 8'd82, 8'd34};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd193, 8'd82, 8'd39};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd167, 8'd63, 8'd24};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd171, 8'd65, 8'd25};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd188, 8'd77, 8'd34};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd191, 8'd74, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd193, 8'd81, 8'd41};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd176, 8'd69, 8'd33};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd127, 8'd27, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd165, 8'd65, 8'd33};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd187, 8'd80, 8'd44};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd187, 8'd75, 8'd35};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd192, 8'd75, 8'd31};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd181, 8'd76, 8'd31};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd167, 8'd58, 8'd15};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd171, 8'd58, 8'd16};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd182, 8'd66, 8'd25};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd178, 8'd62, 8'd21};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd174, 8'd61, 8'd19};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd172, 8'd63, 8'd20};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd165, 8'd60, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd182, 8'd76, 8'd36};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd167, 8'd63, 8'd24};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd163, 8'd69, 8'd35};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd137, 8'd60, 8'd40};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd73, 8'd13, 8'd3};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd80, 8'd23, 8'd14};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd143, 8'd76, 8'd57};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd151, 8'd70, 8'd41};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd133, 8'd33, 8'd9};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd135, 8'd45, 8'd11};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd123, 8'd40, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd139, 8'd52, 8'd9};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd148, 8'd51, 8'd16};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd144, 8'd49, 8'd21};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd107, 8'd23, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd90, 8'd19, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd124, 8'd44, 8'd17};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd146, 8'd63, 8'd33};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd136, 8'd50, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd143, 8'd51, 8'd14};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd136, 8'd42, 8'd4};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd150, 8'd56, 8'd18};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd22};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd138, 8'd46, 8'd9};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd115, 8'd40, 8'd1};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd147, 8'd122, 8'd117};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd169, 8'd185, 8'd200};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd159, 8'd182, 8'd188};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd139, 8'd167, 8'd171};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd133, 8'd170, 8'd186};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd130, 8'd160, 8'd171};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd185, 8'd191, 8'd189};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd165, 8'd105, 8'd68};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd161, 8'd99, 8'd52};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd146, 8'd77, 8'd20};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd139, 8'd61, 8'd0};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd141, 8'd51, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd139, 8'd34, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd154, 8'd39, 8'd12};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd192, 8'd70, 8'd55};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd237, 8'd103, 8'd114};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd199, 8'd71, 8'd70};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd187, 8'd55, 8'd50};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd185, 8'd41, 8'd41};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd165, 8'd3, 8'd16};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd177, 8'd11, 8'd23};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd161, 8'd8, 8'd2};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd147, 8'd9, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd157, 8'd5, 8'd2};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd159, 8'd5, 8'd3};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd163, 8'd8, 8'd6};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd173, 8'd13, 8'd13};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd188, 8'd22, 8'd24};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd205, 8'd35, 8'd38};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd219, 8'd46, 8'd50};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd228, 8'd53, 8'd58};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd236, 8'd49, 8'd60};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd242, 8'd49, 8'd54};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd242, 8'd60, 8'd57};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd229, 8'd68, 8'd58};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd234, 8'd67, 8'd59};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd230, 8'd61, 8'd38};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd226, 8'd107, 8'd39};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd100};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd251, 8'd203, 8'd77};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd250, 8'd193, 8'd41};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd228, 8'd141, 8'd44};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd156, 8'd37, 8'd5};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd171, 8'd40, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd180, 8'd43, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd196, 8'd58, 8'd9};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd210, 8'd74, 8'd14};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd212, 8'd100, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd221, 8'd110, 8'd3};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd232, 8'd120, 8'd10};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd237, 8'd125, 8'd13};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd236, 8'd125, 8'd10};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd236, 8'd121, 8'd12};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd236, 8'd121, 8'd14};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd237, 8'd122, 8'd16};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd244, 8'd111, 8'd8};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd247, 8'd115, 8'd14};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd252, 8'd120, 8'd20};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd253, 8'd123, 8'd25};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd250, 8'd123, 8'd26};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd242, 8'd118, 8'd22};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd235, 8'd110, 8'd17};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd230, 8'd107, 8'd14};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd226, 8'd127, 8'd23};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd232, 8'd126, 8'd6};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd242, 8'd125, 8'd0};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd254, 8'd130, 8'd0};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd255, 8'd139, 8'd0};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd254, 8'd148, 8'd4};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd241, 8'd151, 8'd29};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd229, 8'd150, 8'd45};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd227, 8'd193, 8'd85};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd239, 8'd212, 8'd125};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd252, 8'd236, 8'd184};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd97: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd211};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd250, 8'd223, 8'd168};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd240, 8'd193, 8'd113};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd234, 8'd167, 8'd63};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd236, 8'd152, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd240, 8'd146, 8'd14};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd247, 8'd134, 8'd6};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd249, 8'd136, 8'd6};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd251, 8'd140, 8'd7};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd253, 8'd142, 8'd9};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd253, 8'd141, 8'd15};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd250, 8'd137, 8'd19};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd246, 8'd131, 8'd22};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd244, 8'd128, 8'd25};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd253, 8'd139, 8'd15};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd252, 8'd136, 8'd17};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd250, 8'd130, 8'd18};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd249, 8'd126, 8'd20};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd248, 8'd127, 8'd22};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd247, 8'd131, 8'd20};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd246, 8'd137, 8'd20};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd247, 8'd141, 8'd21};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd245, 8'd145, 8'd23};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd240, 8'd141, 8'd22};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd231, 8'd134, 8'd21};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd219, 8'd120, 8'd16};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd104, 8'd9};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd199, 8'd84, 8'd1};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd192, 8'd68, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd189, 8'd58, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd193, 8'd40, 8'd8};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd198, 8'd83, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd48};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd244, 8'd225, 8'd45};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd241, 8'd221, 8'd72};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd240, 8'd168, 8'd83};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd225, 8'd74, 8'd45};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd64, 8'd67};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd240, 8'd62, 8'd62};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd242, 8'd64, 8'd64};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd242, 8'd66, 8'd66};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd240, 8'd64, 8'd64};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd230, 8'd56, 8'd55};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd213, 8'd39, 8'd38};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd193, 8'd21, 8'd19};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd181, 8'd9, 8'd7};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd180, 8'd8, 8'd8};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd176, 8'd6, 8'd6};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd172, 8'd4, 8'd3};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd167, 8'd3, 8'd1};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd166, 8'd7, 8'd3};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd168, 8'd13, 8'd8};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd173, 8'd20, 8'd14};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd176, 8'd25, 8'd18};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd217, 8'd61, 8'd74};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd226, 8'd91, 8'd87};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd229, 8'd117, 8'd95};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd200, 8'd95, 8'd73};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd153, 8'd43, 8'd26};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd149, 8'd38, 8'd18};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd164, 8'd60, 8'd23};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd136, 8'd42, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd130, 8'd50, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd155, 8'd59, 8'd21};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd175, 8'd76, 8'd34};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd169, 8'd90, 8'd21};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd126, 8'd80, 8'd18};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd110, 8'd93, 8'd75};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd168, 8'd173};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd180, 8'd192, 8'd192};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd198, 8'd200, 8'd212};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd186, 8'd199, 8'd205};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd149, 8'd158, 8'd153};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd137, 8'd116, 8'd97};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd115, 8'd51, 8'd16};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd135, 8'd39, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd170, 8'd75, 8'd31};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd146, 8'd61, 8'd20};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd161, 8'd59, 8'd11};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd12};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd158, 8'd62, 8'd22};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd177, 8'd74, 8'd33};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd35};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd186, 8'd78, 8'd40};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd146, 8'd54, 8'd29};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd97, 8'd19, 8'd7};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd153, 8'd68, 8'd47};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd186, 8'd88, 8'd53};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd175, 8'd60, 8'd15};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd198, 8'd80, 8'd32};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd192, 8'd81, 8'd38};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd167, 8'd63, 8'd24};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd170, 8'd64, 8'd24};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd187, 8'd76, 8'd33};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd192, 8'd75, 8'd31};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd193, 8'd81, 8'd41};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd176, 8'd69, 8'd33};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd129, 8'd29, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd163, 8'd63, 8'd31};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd187, 8'd80, 8'd44};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd187, 8'd75, 8'd35};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd191, 8'd74, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd182, 8'd77, 8'd32};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd168, 8'd59, 8'd16};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd173, 8'd60, 8'd18};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd184, 8'd68, 8'd27};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd180, 8'd64, 8'd23};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd176, 8'd63, 8'd21};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd175, 8'd66, 8'd23};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd168, 8'd63, 8'd18};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd184, 8'd77, 8'd35};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd167, 8'd61, 8'd19};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd151, 8'd53, 8'd18};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd138, 8'd58, 8'd35};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd99, 8'd37, 8'd26};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd88, 8'd30, 8'd19};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd131, 8'd60, 8'd40};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd151, 8'd68, 8'd36};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd134, 8'd34, 8'd10};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd136, 8'd45, 8'd14};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd123, 8'd40, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd138, 8'd50, 8'd10};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd148, 8'd51, 8'd16};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd143, 8'd48, 8'd20};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd106, 8'd21, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd90, 8'd19, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd124, 8'd44, 8'd17};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd147, 8'd64, 8'd34};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd136, 8'd50, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd143, 8'd51, 8'd14};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd136, 8'd42, 8'd4};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd149, 8'd55, 8'd17};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd22};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd137, 8'd45, 8'd8};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd113, 8'd37, 8'd1};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd154, 8'd131, 8'd125};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd168, 8'd186, 8'd200};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd155, 8'd178, 8'd184};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd124, 8'd152, 8'd156};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd125, 8'd163, 8'd176};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd122, 8'd150, 8'd162};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd175, 8'd180, 8'd176};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd157, 8'd96, 8'd33};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd149, 8'd81, 8'd18};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd147, 8'd73, 8'd10};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd146, 8'd59, 8'd5};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd139, 8'd41, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd153, 8'd42, 8'd12};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd194, 8'd72, 8'd57};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd227, 8'd100, 8'd93};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd216, 8'd88, 8'd75};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd207, 8'd85, 8'd64};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd198, 8'd74, 8'd50};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd153, 8'd12, 8'd2};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd166, 8'd6, 8'd14};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd178, 8'd12, 8'd24};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd163, 8'd8, 8'd6};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd156, 8'd15, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd159, 8'd1, 8'd0};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd164, 8'd6, 8'd5};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd175, 8'd15, 8'd15};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd190, 8'd27, 8'd28};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd205, 8'd39, 8'd41};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd218, 8'd49, 8'd52};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd228, 8'd58, 8'd61};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd233, 8'd63, 8'd66};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd239, 8'd60, 8'd66};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd246, 8'd55, 8'd60};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd246, 8'd61, 8'd59};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd236, 8'd65, 8'd58};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd238, 8'd63, 8'd58};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd234, 8'd59, 8'd38};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd228, 8'd109, 8'd43};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd105};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd237, 8'd209, 8'd40};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd243, 8'd200, 8'd10};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd232, 8'd150, 8'd22};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd168, 8'd48, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd186, 8'd50, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd194, 8'd55, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd204, 8'd68, 8'd10};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd216, 8'd85, 8'd17};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd223, 8'd112, 8'd5};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd233, 8'd121, 8'd11};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd244, 8'd133, 8'd17};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd253, 8'd140, 8'd18};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd254, 8'd140, 8'd16};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd254, 8'd139, 8'd14};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd139, 8'd16};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd20};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd248, 8'd138, 8'd23};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd246, 8'd137, 8'd20};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd244, 8'd133, 8'd17};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd244, 8'd129, 8'd12};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd245, 8'd129, 8'd10};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd248, 8'd129, 8'd9};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd251, 8'd131, 8'd9};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd254, 8'd131, 8'd10};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd247, 8'd140, 8'd10};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd251, 8'd144, 8'd6};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd252, 8'd146, 8'd0};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd246, 8'd146, 8'd0};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd237, 8'd150, 8'd11};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd234, 8'd162, 8'd44};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd238, 8'd182, 8'd87};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd245, 8'd198, 8'd118};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd172};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd195};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd255, 8'd249, 8'd226};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd98: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd224};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd251, 8'd219, 8'd178};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd243, 8'd204, 8'd125};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd237, 8'd194, 8'd90};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd23};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd241, 8'd153, 8'd17};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd242, 8'd149, 8'd9};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd245, 8'd146, 8'd3};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd251, 8'd145, 8'd1};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd255, 8'd145, 8'd4};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd148, 8'd10};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd13};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd247, 8'd141, 8'd3};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd246, 8'd140, 8'd5};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd246, 8'd137, 8'd8};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd248, 8'd138, 8'd13};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd250, 8'd142, 8'd16};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd253, 8'd150, 8'd22};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd25};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd26};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd25};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd26};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd244, 8'd156, 8'd23};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd232, 8'd138, 8'd22};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd118, 8'd16};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd205, 8'd97, 8'd9};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd195, 8'd79, 8'd4};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd189, 8'd67, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd191, 8'd47, 8'd12};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd203, 8'd92, 8'd2};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd53};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd248, 8'd222, 8'd49};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd248, 8'd220, 8'd77};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd242, 8'd164, 8'd82};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd225, 8'd71, 8'd45};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd63, 8'd66};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd242, 8'd64, 8'd64};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd241, 8'd63, 8'd63};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd241, 8'd65, 8'd65};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd244, 8'd68, 8'd68};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd243, 8'd69, 8'd68};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd58, 8'd57};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd212, 8'd40, 8'd38};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd196, 8'd24, 8'd22};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd188, 8'd12, 8'd14};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd186, 8'd12, 8'd13};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd181, 8'd11, 8'd11};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd176, 8'd11, 8'd9};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd170, 8'd11, 8'd7};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd165, 8'd10, 8'd5};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd161, 8'd10, 8'd3};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd158, 8'd9, 8'd2};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd186, 8'd28, 8'd42};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd200, 8'd61, 8'd56};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd222, 8'd106, 8'd83};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd217, 8'd107, 8'd84};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd191, 8'd73, 8'd59};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd160, 8'd38, 8'd27};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd142, 8'd25, 8'd5};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd149, 8'd42, 8'd8};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd128, 8'd49, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd148, 8'd53, 8'd9};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd171, 8'd69, 8'd21};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd181, 8'd99, 8'd25};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd147, 8'd98, 8'd31};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd106, 8'd86, 8'd61};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd169, 8'd168};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd177, 8'd190, 8'd183};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd194, 8'd197, 8'd206};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd189, 8'd202, 8'd208};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd147, 8'd159, 8'd155};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd142, 8'd125, 8'd107};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd112, 8'd49, 8'd16};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd137, 8'd44, 8'd3};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd169, 8'd72, 8'd29};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd149, 8'd61, 8'd21};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd168, 8'd62, 8'd20};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd156, 8'd57, 8'd18};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd151, 8'd54, 8'd19};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd172, 8'd70, 8'd32};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd191, 8'd85, 8'd43};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd166, 8'd66, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd117, 8'd33, 8'd9};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd85, 8'd17, 8'd6};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd150, 8'd65, 8'd44};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd189, 8'd91, 8'd56};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd176, 8'd61, 8'd16};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd195, 8'd77, 8'd29};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd192, 8'd81, 8'd38};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd168, 8'd64, 8'd25};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd170, 8'd64, 8'd24};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd187, 8'd76, 8'd33};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd192, 8'd75, 8'd31};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd192, 8'd80, 8'd40};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd175, 8'd68, 8'd32};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd132, 8'd32, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd160, 8'd60, 8'd28};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd188, 8'd81, 8'd45};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd188, 8'd76, 8'd36};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd191, 8'd74, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd184, 8'd79, 8'd34};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd170, 8'd61, 8'd18};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd175, 8'd62, 8'd20};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd187, 8'd71, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd184, 8'd68, 8'd27};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd180, 8'd67, 8'd25};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd179, 8'd70, 8'd27};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd172, 8'd67, 8'd22};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd184, 8'd72, 8'd26};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd175, 8'd64, 8'd19};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd146, 8'd44, 8'd4};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd132, 8'd48, 8'd22};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd117, 8'd50, 8'd34};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd106, 8'd43, 8'd28};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd128, 8'd54, 8'd29};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd147, 8'd58, 8'd24};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd135, 8'd37, 8'd12};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd136, 8'd47, 8'd15};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd122, 8'd40, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd135, 8'd50, 8'd9};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd144, 8'd50, 8'd14};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd142, 8'd47, 8'd19};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd104, 8'd22, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd87, 8'd19, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd125, 8'd45, 8'd18};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd148, 8'd65, 8'd35};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd136, 8'd50, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd143, 8'd51, 8'd14};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd136, 8'd42, 8'd4};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd148, 8'd54, 8'd16};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd149, 8'd57, 8'd20};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd136, 8'd44, 8'd7};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd114, 8'd41, 8'd6};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd169, 8'd148, 8'd143};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd172, 8'd191, 8'd205};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd155, 8'd178, 8'd186};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd111, 8'd136, 8'd140};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd124, 8'd160, 8'd174};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd121, 8'd148, 8'd159};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd170, 8'd172, 8'd169};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd183, 8'd113, 8'd27};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd166, 8'd90, 8'd14};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd162, 8'd76, 8'd15};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd153, 8'd56, 8'd13};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd143, 8'd33, 8'd6};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd176, 8'd55, 8'd38};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd219, 8'd91, 8'd80};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd226, 8'd93, 8'd84};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd212, 8'd96, 8'd47};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd231, 8'd120, 8'd65};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd228, 8'd114, 8'd62};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd133, 8'd2, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd169, 8'd15, 8'd13};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd183, 8'd17, 8'd29};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd171, 8'd10, 8'd15};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd172, 8'd23, 8'd16};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd177, 8'd11, 8'd11};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd185, 8'd19, 8'd19};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd198, 8'd32, 8'd32};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd212, 8'd46, 8'd46};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd223, 8'd57, 8'd57};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd230, 8'd64, 8'd64};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd232, 8'd66, 8'd66};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd233, 8'd67, 8'd67};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd241, 8'd75, 8'd75};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd250, 8'd64, 8'd65};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd252, 8'd63, 8'd61};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd242, 8'd58, 8'd56};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd245, 8'd55, 8'd55};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd236, 8'd55, 8'd38};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd228, 8'd110, 8'd46};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd110};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd242, 8'd232, 8'd46};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd253, 8'd222, 8'd17};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd248, 8'd171, 8'd33};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd190, 8'd65, 8'd7};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd208, 8'd63, 8'd6};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd208, 8'd65, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd212, 8'd75, 8'd21};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd216, 8'd91, 8'd25};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd223, 8'd130, 8'd26};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd232, 8'd140, 8'd31};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd246, 8'd153, 8'd34};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd254, 8'd160, 8'd34};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd26};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd27};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd242, 8'd152, 8'd14};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd243, 8'd153, 8'd15};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd246, 8'd153, 8'd13};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd252, 8'd155, 8'd14};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd13};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd15};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd16};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd16};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd6};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd250, 8'd153, 8'd10};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd240, 8'd159, 8'd24};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd235, 8'd173, 8'd52};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd237, 8'd193, 8'd94};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd244, 8'd216, 8'd142};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd252, 8'd235, 8'd181};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd204};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd99: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd216};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd192};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd251, 8'd200, 8'd109};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd245, 8'd191, 8'd95};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd237, 8'd174, 8'd68};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd233, 8'd161, 8'd41};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd236, 8'd152, 8'd20};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd248, 8'd151, 8'd10};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd6};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd6};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd250, 8'd163, 8'd24};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd252, 8'd164, 8'd28};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd34};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd34};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd250, 8'd166, 8'd31};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd26};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd23};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd23};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd251, 8'd164, 8'd23};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd243, 8'd151, 8'd24};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd231, 8'd133, 8'd24};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd217, 8'd111, 8'd23};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd202, 8'd90, 8'd18};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd190, 8'd71, 8'd13};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd183, 8'd61, 8'd10};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd184, 8'd50, 8'd12};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd206, 8'd98, 8'd8};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd49};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd249, 8'd211, 8'd48};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd252, 8'd209, 8'd78};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd238, 8'd150, 8'd76};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd218, 8'd62, 8'd39};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd255, 8'd56, 8'd58};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd248, 8'd70, 8'd70};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd246, 8'd68, 8'd68};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd243, 8'd67, 8'd67};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd244, 8'd68, 8'd68};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd242, 8'd68, 8'd67};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd237, 8'd63, 8'd62};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd227, 8'd55, 8'd53};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd219, 8'd47, 8'd45};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd197, 8'd17, 8'd20};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd194, 8'd15, 8'd18};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd189, 8'd15, 8'd16};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd181, 8'd13, 8'd12};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd174, 8'd12, 8'd9};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd166, 8'd11, 8'd6};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd163, 8'd12, 8'd5};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd159, 8'd12, 8'd4};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd164, 8'd7, 8'd14};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd180, 8'd42, 8'd29};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd204, 8'd87, 8'd54};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd208, 8'd95, 8'd63};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd216, 8'd95, 8'd78};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd199, 8'd70, 8'd64};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd150, 8'd23, 8'd14};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd148, 8'd28, 8'd11};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd130, 8'd50, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd141, 8'd43, 8'd6};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd160, 8'd54, 8'd12};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd179, 8'd90, 8'd24};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd162, 8'd106, 8'd47};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd158, 8'd132, 8'd115};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd184, 8'd183, 8'd189};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd173, 8'd185, 8'd185};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd189, 8'd194, 8'd200};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd188, 8'd206, 8'd210};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd146, 8'd162, 8'd161};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd148, 8'd135, 8'd119};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd109, 8'd50, 8'd20};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd141, 8'd47, 8'd9};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd168, 8'd69, 8'd27};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd153, 8'd61, 8'd20};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd171, 8'd63, 8'd24};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd162, 8'd59, 8'd24};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd147, 8'd50, 8'd17};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd166, 8'd66, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd190, 8'd88, 8'd48};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd154, 8'd57, 8'd22};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd94, 8'd16, 8'd0};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd77, 8'd15, 8'd4};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd147, 8'd62, 8'd41};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd192, 8'd94, 8'd59};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd176, 8'd61, 8'd16};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd191, 8'd73, 8'd25};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd192, 8'd81, 8'd38};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd170, 8'd66, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd23};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd186, 8'd75, 8'd32};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd193, 8'd76, 8'd32};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd191, 8'd79, 8'd39};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd173, 8'd66, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd136, 8'd36, 8'd4};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd156, 8'd56, 8'd24};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd190, 8'd83, 8'd47};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd189, 8'd77, 8'd37};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd190, 8'd73, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd185, 8'd80, 8'd35};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd172, 8'd63, 8'd20};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd177, 8'd64, 8'd22};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd189, 8'd73, 8'd32};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd187, 8'd71, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd184, 8'd71, 8'd29};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd183, 8'd74, 8'd31};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd177, 8'd72, 8'd27};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd181, 8'd66, 8'd19};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd181, 8'd66, 8'd19};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd155, 8'd49, 8'd7};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd126, 8'd39, 8'd11};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd107, 8'd36, 8'd18};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd117, 8'd50, 8'd33};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd145, 8'd68, 8'd42};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd143, 8'd51, 8'd14};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd137, 8'd41, 8'd17};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd136, 8'd49, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd123, 8'd41, 8'd3};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd134, 8'd49, 8'd10};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd142, 8'd48, 8'd14};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd140, 8'd46, 8'd20};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd102, 8'd21, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd87, 8'd19, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd126, 8'd46, 8'd19};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd149, 8'd66, 8'd36};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd137, 8'd51, 8'd18};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd143, 8'd51, 8'd14};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd135, 8'd41, 8'd3};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd147, 8'd53, 8'd15};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd147, 8'd55, 8'd18};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd134, 8'd42, 8'd5};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd116, 8'd50, 8'd15};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd185, 8'd167, 8'd163};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd176, 8'd198, 8'd212};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd156, 8'd181, 8'd188};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd104, 8'd129, 8'd133};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd131, 8'd165, 8'd177};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd133, 8'd155, 8'd166};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd178, 8'd175, 8'd170};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd181, 8'd99, 8'd15};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd165, 8'd77, 8'd6};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd145, 8'd49, 8'd1};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd137, 8'd29, 8'd1};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd148, 8'd31, 8'd13};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd180, 8'd55, 8'd35};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd197, 8'd69, 8'd40};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd193, 8'd63, 8'd27};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd237, 8'd133, 8'd44};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd68};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd255, 8'd157, 8'd75};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd158, 8'd36, 8'd0};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd176, 8'd26, 8'd12};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd193, 8'd28, 8'd35};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd184, 8'd18, 8'd28};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd190, 8'd34, 8'd35};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd210, 8'd37, 8'd39};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd215, 8'd42, 8'd44};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd221, 8'd51, 8'd52};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd229, 8'd59, 8'd60};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd233, 8'd65, 8'd65};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd233, 8'd67, 8'd67};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd233, 8'd67, 8'd67};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd231, 8'd67, 8'd66};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd241, 8'd84, 8'd79};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd250, 8'd68, 8'd65};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd254, 8'd58, 8'd59};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd244, 8'd50, 8'd51};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd248, 8'd45, 8'd49};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd237, 8'd47, 8'd35};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd227, 8'd107, 8'd46};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd112};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd242, 8'd239, 8'd72};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd254, 8'd226, 8'd39};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd249, 8'd170, 8'd49};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd191, 8'd63, 8'd18};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd207, 8'd61, 8'd12};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd206, 8'd64, 8'd2};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd207, 8'd78, 8'd21};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd209, 8'd95, 8'd24};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd211, 8'd140, 8'd32};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd219, 8'd149, 8'd35};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd231, 8'd161, 8'd37};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd238, 8'd168, 8'd34};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd241, 8'd168, 8'd27};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd241, 8'd166, 8'd21};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd243, 8'd167, 8'd21};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd245, 8'd169, 8'd21};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd14};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd15};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd255, 8'd169, 8'd15};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd17};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd250, 8'd164, 8'd19};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd247, 8'd162, 8'd20};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd245, 8'd159, 8'd20};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd242, 8'd159, 8'd21};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd250, 8'd172, 8'd48};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd244, 8'd178, 8'd66};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd238, 8'd194, 8'd99};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd240, 8'd218, 8'd145};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd249, 8'd241, 8'd192};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd100: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd253, 8'd235, 8'd211};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd254, 8'd231, 8'd199};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd254, 8'd223, 8'd177};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd251, 8'd210, 8'd144};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd246, 8'd195, 8'd106};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd66};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd232, 8'd163, 8'd34};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd227, 8'd154, 8'd16};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd240, 8'd154, 8'd19};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd244, 8'd156, 8'd20};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd252, 8'd161, 8'd21};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd22};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd22};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd19};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd252, 8'd168, 8'd18};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd247, 8'd167, 8'd16};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd252, 8'd169, 8'd15};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd249, 8'd163, 8'd16};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd243, 8'd151, 8'd18};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd233, 8'd132, 8'd18};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd219, 8'd110, 8'd15};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd203, 8'd90, 8'd12};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd191, 8'd73, 8'd9};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd183, 8'd64, 8'd6};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd173, 8'd50, 8'd8};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd201, 8'd100, 8'd10};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd44};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd245, 8'd196, 8'd41};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd251, 8'd195, 8'd74};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd231, 8'd132, 8'd65};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd208, 8'd48, 8'd26};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd250, 8'd44, 8'd46};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd241, 8'd63, 8'd63};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd247, 8'd69, 8'd69};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd250, 8'd74, 8'd74};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd249, 8'd73, 8'd73};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd242, 8'd68, 8'd67};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd235, 8'd61, 8'd60};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd230, 8'd58, 8'd56};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd229, 8'd57, 8'd55};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd213, 8'd34, 8'd37};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd206, 8'd30, 8'd32};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd197, 8'd23, 8'd24};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd185, 8'd17, 8'd16};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd177, 8'd13, 8'd11};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd171, 8'd14, 8'd9};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd168, 8'd15, 8'd9};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd168, 8'd17, 8'd10};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd157, 8'd9, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd189, 8'd60, 8'd28};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd237, 8'd127, 8'd74};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd212, 8'd106, 8'd54};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd194, 8'd75, 8'd41};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd228, 8'd98, 8'd84};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd200, 8'd72, 8'd63};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd136, 8'd12, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd121, 8'd39, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd134, 8'd32, 8'd9};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd152, 8'd41, 8'd13};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd163, 8'd66, 8'd15};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd152, 8'd88, 8'd44};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd213, 8'd182, 8'd179};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd198, 8'd193, 8'd213};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd172, 8'd182, 8'd194};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd186, 8'd191, 8'd197};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd187, 8'd206, 8'd210};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd148, 8'd168, 8'd167};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd151, 8'd141, 8'd129};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd110, 8'd54, 8'd27};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd140, 8'd48, 8'd11};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd169, 8'd68, 8'd26};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd156, 8'd60, 8'd18};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd170, 8'd62, 8'd23};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd167, 8'd64, 8'd29};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd149, 8'd52, 8'd19};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd162, 8'd62, 8'd26};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd189, 8'd87, 8'd47};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd155, 8'd58, 8'd23};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd92, 8'd14, 8'd0};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd74, 8'd12, 8'd1};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd143, 8'd58, 8'd37};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd196, 8'd98, 8'd63};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd177, 8'd62, 8'd17};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd187, 8'd69, 8'd21};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd172, 8'd68, 8'd29};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd168, 8'd62, 8'd22};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd185, 8'd74, 8'd31};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd194, 8'd77, 8'd33};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd190, 8'd78, 8'd38};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd171, 8'd64, 8'd28};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd140, 8'd40, 8'd8};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd152, 8'd52, 8'd20};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd192, 8'd85, 8'd49};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd190, 8'd78, 8'd38};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd189, 8'd72, 8'd28};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd184, 8'd79, 8'd34};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd171, 8'd62, 8'd19};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd177, 8'd64, 8'd22};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd189, 8'd73, 8'd32};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd188, 8'd72, 8'd31};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd186, 8'd73, 8'd31};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd185, 8'd76, 8'd33};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd179, 8'd74, 8'd29};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd185, 8'd69, 8'd20};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd175, 8'd61, 8'd11};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd162, 8'd55, 8'd13};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd131, 8'd42, 8'd12};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd87, 8'd16, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd108, 8'd41, 8'd24};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd161, 8'd81, 8'd54};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd148, 8'd56, 8'd17};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd140, 8'd44, 8'd22};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd138, 8'd51, 8'd23};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd121, 8'd41, 8'd4};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd132, 8'd49, 8'd9};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd139, 8'd46, 8'd13};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd136, 8'd44, 8'd19};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd101, 8'd20, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd86, 8'd19, 8'd2};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd128, 8'd48, 8'd21};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd150, 8'd67, 8'd37};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd137, 8'd51, 8'd18};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd13};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd134, 8'd40, 8'd2};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd145, 8'd51, 8'd13};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd145, 8'd53, 8'd16};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd131, 8'd39, 8'd2};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd117, 8'd54, 8'd19};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd187, 8'd173, 8'd170};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd170, 8'd193, 8'd209};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd148, 8'd173, 8'd180};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd101, 8'd125, 8'd129};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd134, 8'd164, 8'd175};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd142, 8'd160, 8'd170};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd182, 8'd175, 8'd169};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd152, 8'd59, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd144, 8'd48, 8'd0};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd129, 8'd26, 8'd0};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd148, 8'd38, 8'd15};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd187, 8'd71, 8'd46};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd187, 8'd67, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd188, 8'd67, 8'd10};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd225, 8'd104, 8'd35};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd252, 8'd161, 8'd44};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd55};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd70};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd205, 8'd94, 8'd23};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd178, 8'd37, 8'd10};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd203, 8'd39, 8'd40};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd203, 8'd33, 8'd42};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd210, 8'd45, 8'd49};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd56};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd230, 8'd56, 8'd57};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd232, 8'd58, 8'd59};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd234, 8'd62, 8'd62};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd234, 8'd64, 8'd64};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd236, 8'd66, 8'd66};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd236, 8'd68, 8'd67};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd237, 8'd69, 8'd68};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd236, 8'd79, 8'd72};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd245, 8'd62, 8'd58};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd246, 8'd51, 8'd49};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd236, 8'd40, 8'd42};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd240, 8'd35, 8'd40};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd231, 8'd37, 8'd27};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd224, 8'd99, 8'd41};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd108};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd252, 8'd241, 8'd87};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd51};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd250, 8'd176, 8'd55};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd187, 8'd70, 8'd16};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd202, 8'd74, 8'd3};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd202, 8'd81, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd208, 8'd100, 8'd9};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd212, 8'd120, 8'd11};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd229, 8'd150, 8'd19};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd237, 8'd160, 8'd22};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd246, 8'd170, 8'd24};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd252, 8'd175, 8'd21};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd251, 8'd175, 8'd14};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd248, 8'd172, 8'd9};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd248, 8'd172, 8'd8};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd249, 8'd173, 8'd9};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd9};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd12};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd247, 8'd158, 8'd16};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd236, 8'd157, 8'd26};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd231, 8'd162, 8'd43};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd233, 8'd172, 8'd65};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd236, 8'd182, 8'd84};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd239, 8'd190, 8'd95};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd245, 8'd208, 8'd140};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd251, 8'd225, 8'd166};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd203};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd101: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd200};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd250, 8'd224, 8'd163};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd238, 8'd206, 8'd129};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd230, 8'd196, 8'd107};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd244, 8'd163, 8'd48};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd245, 8'd160, 8'd41};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd246, 8'd157, 8'd31};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd248, 8'd156, 8'd23};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd251, 8'd155, 8'd16};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd254, 8'd159, 8'd15};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd16};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd19};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd241, 8'd173, 8'd14};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd239, 8'd166, 8'd12};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd234, 8'd151, 8'd11};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd225, 8'd133, 8'd8};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd210, 8'd112, 8'd3};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd193, 8'd93, 8'd0};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd178, 8'd76, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd170, 8'd68, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd163, 8'd51, 8'd5};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd200, 8'd102, 8'd13};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd252, 8'd176, 8'd39};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd243, 8'd183, 8'd37};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd252, 8'd182, 8'd70};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd223, 8'd114, 8'd55};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd199, 8'd34, 8'd15};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd238, 8'd34, 8'd35};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd44, 8'd44};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd235, 8'd57, 8'd57};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd248, 8'd72, 8'd72};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd253, 8'd77, 8'd77};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd246, 8'd72, 8'd71};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd236, 8'd62, 8'd61};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd228, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd227, 8'd55, 8'd53};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd229, 8'd55, 8'd56};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd221, 8'd49, 8'd49};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd208, 8'd38, 8'd38};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd196, 8'd28, 8'd27};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd185, 8'd20, 8'd18};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd180, 8'd16, 8'd14};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd178, 8'd16, 8'd13};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd176, 8'd17, 8'd13};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd155, 8'd23, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd224, 8'd110, 8'd48};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd80};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd222, 8'd127, 8'd45};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd197, 8'd88, 8'd29};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd203, 8'd80, 8'd47};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd184, 8'd59, 8'd41};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd162, 8'd41, 8'd24};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd117, 8'd34, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd134, 8'd29, 8'd10};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd151, 8'd34, 8'd14};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd151, 8'd48, 8'd3};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd133, 8'd64, 8'd25};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd225, 8'd190, 8'd194};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd198, 8'd190, 8'd214};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd174, 8'd183, 8'd200};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd181, 8'd189, 8'd192};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd185, 8'd206, 8'd209};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd152, 8'd176, 8'd176};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd149, 8'd145, 8'd134};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd115, 8'd61, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd138, 8'd45, 8'd11};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd172, 8'd69, 8'd28};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd157, 8'd58, 8'd16};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd163, 8'd57, 8'd15};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd171, 8'd72, 8'd33};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd157, 8'd60, 8'd25};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd161, 8'd59, 8'd21};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd189, 8'd83, 8'd41};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd168, 8'd68, 8'd32};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd110, 8'd26, 8'd2};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd77, 8'd9, 8'd0};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd140, 8'd55, 8'd34};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd199, 8'd101, 8'd66};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd178, 8'd63, 8'd18};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd183, 8'd65, 8'd17};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd174, 8'd70, 8'd31};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd167, 8'd61, 8'd21};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd184, 8'd73, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd194, 8'd77, 8'd33};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd190, 8'd78, 8'd38};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd170, 8'd63, 8'd27};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd144, 8'd44, 8'd12};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd148, 8'd48, 8'd16};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd193, 8'd86, 8'd50};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd191, 8'd79, 8'd39};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd189, 8'd72, 8'd28};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd182, 8'd77, 8'd32};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd169, 8'd60, 8'd17};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd175, 8'd62, 8'd20};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd188, 8'd72, 8'd31};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd187, 8'd71, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd186, 8'd73, 8'd31};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd186, 8'd77, 8'd34};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd180, 8'd75, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd186, 8'd71, 8'd24};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd166, 8'd51, 8'd4};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd160, 8'd54, 8'd12};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd137, 8'd50, 8'd22};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd83, 8'd12, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd97, 8'd30, 8'd13};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd159, 8'd82, 8'd56};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd159, 8'd67, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd142, 8'd47, 8'd25};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd140, 8'd55, 8'd26};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd120, 8'd42, 8'd4};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd130, 8'd48, 8'd10};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd136, 8'd46, 8'd12};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd134, 8'd42, 8'd17};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd98, 8'd20, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd85, 8'd20, 8'd2};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd129, 8'd49, 8'd22};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd151, 8'd68, 8'd38};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd138, 8'd52, 8'd19};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd13};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd133, 8'd39, 8'd1};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd144, 8'd50, 8'd12};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd143, 8'd51, 8'd14};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd129, 8'd37, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd121, 8'd62, 8'd28};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd182, 8'd172, 8'd170};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd156, 8'd184, 8'd198};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd133, 8'd160, 8'd167};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd98, 8'd122, 8'd126};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd127, 8'd155, 8'd167};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd144, 8'd158, 8'd167};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd177, 8'd164, 8'd158};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd140, 8'd43, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd144, 8'd46, 8'd7};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd147, 8'd44, 8'd13};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd189, 8'd81, 8'd52};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd222, 8'd112, 8'd75};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd184, 8'd73, 8'd20};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd185, 8'd74, 8'd3};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd74};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd245, 8'd162, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd241, 8'd164, 8'd32};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd247, 8'd168, 8'd49};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd241, 8'd139, 8'd57};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd190, 8'd52, 8'd15};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd210, 8'd47, 8'd42};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd218, 8'd45, 8'd47};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd225, 8'd53, 8'd53};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd227, 8'd53, 8'd52};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd228, 8'd54, 8'd53};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd230, 8'd56, 8'd55};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd232, 8'd58, 8'd57};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd235, 8'd61, 8'd60};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd238, 8'd64, 8'd63};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd240, 8'd66, 8'd65};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd241, 8'd67, 8'd66};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd227, 8'd60, 8'd54};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd233, 8'd46, 8'd41};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd232, 8'd39, 8'd34};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd221, 8'd31, 8'd31};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd227, 8'd26, 8'd32};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd221, 8'd27, 8'd18};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd219, 8'd85, 8'd32};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd100};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd77};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd40};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd252, 8'd185, 8'd45};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd181, 8'd86, 8'd6};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd189, 8'd89, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd188, 8'd96, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd191, 8'd108, 8'd0};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd194, 8'd125, 8'd0};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd239, 8'd139, 8'd0};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd245, 8'd149, 8'd3};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd11};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd11};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd11};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd251, 8'd166, 8'd11};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd250, 8'd167, 8'd13};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd250, 8'd169, 8'd17};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd240, 8'd159, 8'd41};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd241, 8'd163, 8'd52};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd241, 8'd173, 8'd72};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd244, 8'd188, 8'd101};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd249, 8'd205, 8'd132};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd254, 8'd224, 8'd164};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd189};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd203};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd102: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd176};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd162};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd139};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd251, 8'd199, 8'd115};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd244, 8'd188, 8'd93};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd239, 8'd180, 8'd80};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd237, 8'd175, 8'd72};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd235, 8'd173, 8'd70};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd228, 8'd178, 8'd53};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd226, 8'd170, 8'd51};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd221, 8'd155, 8'd45};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd209, 8'd133, 8'd35};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd193, 8'd112, 8'd23};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd173, 8'd90, 8'd10};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd156, 8'd74, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd144, 8'd64, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd158, 8'd53, 8'd5};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd201, 8'd107, 8'd17};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd249, 8'd170, 8'd39};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd243, 8'd174, 8'd35};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd254, 8'd175, 8'd70};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd221, 8'd104, 8'd50};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd193, 8'd26, 8'd10};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd232, 8'd28, 8'd29};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd210, 8'd32, 8'd32};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd220, 8'd42, 8'd42};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd232, 8'd56, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd242, 8'd66, 8'd66};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd244, 8'd70, 8'd69};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd240, 8'd66, 8'd65};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd232, 8'd60, 8'd58};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd228, 8'd56, 8'd54};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd224, 8'd59, 8'd57};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd221, 8'd56, 8'd54};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd218, 8'd50, 8'd49};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd211, 8'd43, 8'd42};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd203, 8'd35, 8'd34};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd197, 8'd29, 8'd28};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd193, 8'd23, 8'd23};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd191, 8'd21, 8'd21};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd174, 8'd59, 8'd0};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd246, 8'd148, 8'd57};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd246, 8'd166, 8'd53};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd232, 8'd152, 8'd39};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd236, 8'd140, 8'd54};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd185, 8'd74, 8'd21};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd155, 8'd38, 8'd5};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd192, 8'd78, 8'd52};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd144, 8'd62, 8'd14};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd145, 8'd41, 8'd16};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd149, 8'd29, 8'd4};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd151, 8'd45, 8'd0};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd136, 8'd63, 8'd20};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd207, 8'd169, 8'd166};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd192, 8'd185, 8'd203};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd171, 8'd181, 8'd191};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd179, 8'd187, 8'd189};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd181, 8'd205, 8'd207};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd158, 8'd184, 8'd185};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd148, 8'd145, 8'd138};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd119, 8'd68, 8'd47};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd133, 8'd43, 8'd9};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd174, 8'd71, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd160, 8'd57, 8'd16};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd153, 8'd51, 8'd3};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd174, 8'd77, 8'd34};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd166, 8'd70, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd160, 8'd57, 8'd16};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd188, 8'd77, 8'd32};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd189, 8'd81, 8'd43};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd135, 8'd43, 8'd18};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd85, 8'd7, 8'd0};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd137, 8'd52, 8'd31};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd202, 8'd104, 8'd69};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd179, 8'd64, 8'd19};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd180, 8'd62, 8'd14};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd175, 8'd71, 8'd32};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd166, 8'd60, 8'd20};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd183, 8'd72, 8'd29};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd195, 8'd78, 8'd34};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd189, 8'd77, 8'd37};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd169, 8'd62, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd148, 8'd48, 8'd16};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd144, 8'd44, 8'd12};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd194, 8'd87, 8'd51};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd191, 8'd79, 8'd39};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd188, 8'd71, 8'd27};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd179, 8'd74, 8'd29};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd166, 8'd57, 8'd14};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd172, 8'd59, 8'd17};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd186, 8'd70, 8'd29};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd186, 8'd70, 8'd29};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd185, 8'd72, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd185, 8'd76, 8'd33};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd180, 8'd75, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd173, 8'd61, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd168, 8'd57, 8'd11};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd158, 8'd54, 8'd15};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd133, 8'd47, 8'd20};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd89, 8'd22, 8'd6};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd99, 8'd36, 8'd21};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd151, 8'd75, 8'd51};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd155, 8'd67, 8'd31};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd145, 8'd50, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd141, 8'd55, 8'd28};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd121, 8'd43, 8'd7};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd129, 8'd47, 8'd9};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd134, 8'd43, 8'd12};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd132, 8'd42, 8'd18};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd98, 8'd19, 8'd2};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd85, 8'd19, 8'd3};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd130, 8'd50, 8'd23};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd151, 8'd68, 8'd38};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd138, 8'd52, 8'd19};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd13};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd133, 8'd39, 8'd1};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd143, 8'd49, 8'd11};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd13};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd128, 8'd36, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd137, 8'd83, 8'd49};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd183, 8'd178, 8'd175};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd153, 8'd182, 8'd198};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd126, 8'd153, 8'd162};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd103, 8'd127, 8'd131};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd120, 8'd147, 8'd158};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd145, 8'd155, 8'd164};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd169, 8'd154, 8'd147};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd138, 8'd46, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd153, 8'd61, 8'd14};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd168, 8'd73, 8'd27};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd191, 8'd93, 8'd48};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd193, 8'd93, 8'd44};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd152, 8'd51, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd158, 8'd56, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd225, 8'd122, 8'd55};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd235, 8'd159, 8'd22};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd237, 8'd168, 8'd31};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd238, 8'd164, 8'd41};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd74};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd210, 8'd77, 8'd34};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd213, 8'd49, 8'd37};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd223, 8'd48, 8'd45};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd225, 8'd51, 8'd44};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd218, 8'd49, 8'd46};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd221, 8'd52, 8'd49};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd228, 8'd56, 8'd54};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd233, 8'd59, 8'd58};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd237, 8'd59, 8'd59};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd236, 8'd56, 8'd57};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd234, 8'd51, 8'd53};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd231, 8'd48, 8'd50};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd215, 8'd37, 8'd33};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd220, 8'd28, 8'd25};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd216, 8'd27, 8'd21};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd205, 8'd23, 8'd19};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd210, 8'd20, 8'd22};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd212, 8'd18, 8'd9};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd214, 8'd72, 8'd22};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd89};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd254, 8'd204, 8'd47};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd23};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd243, 8'd179, 8'd45};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd173, 8'd94, 8'd25};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd183, 8'd107, 8'd23};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd180, 8'd110, 8'd12};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd183, 8'd118, 8'd26};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd189, 8'd127, 8'd24};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd222, 8'd140, 8'd38};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd229, 8'd150, 8'd47};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd239, 8'd165, 8'd60};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd243, 8'd174, 8'd70};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd241, 8'd179, 8'd78};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd237, 8'd181, 8'd84};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd238, 8'd184, 8'd94};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd238, 8'd188, 8'd103};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd103: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd250, 8'd212, 8'd139};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd247, 8'd202, 8'd134};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd241, 8'd185, 8'd124};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd228, 8'd163, 8'd109};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd208, 8'd137, 8'd91};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd186, 8'd115, 8'd73};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd165, 8'd97, 8'd58};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd153, 8'd88, 8'd50};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd156, 8'd56, 8'd4};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd202, 8'd111, 8'd22};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd251, 8'd170, 8'd39};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd245, 8'd171, 8'd36};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd72};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd221, 8'd101, 8'd49};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd193, 8'd23, 8'd8};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd230, 8'd26, 8'd27};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd209, 8'd31, 8'd31};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd210, 8'd32, 8'd32};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd214, 8'd38, 8'd38};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd237, 8'd63, 8'd62};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd243, 8'd69, 8'd68};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd240, 8'd68, 8'd66};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd235, 8'd63, 8'd61};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd211, 8'd49, 8'd46};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd214, 8'd52, 8'd49};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd217, 8'd53, 8'd51};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd221, 8'd53, 8'd52};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd219, 8'd49, 8'd49};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd215, 8'd43, 8'd43};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd209, 8'd35, 8'd36};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd206, 8'd30, 8'd32};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd210, 8'd106, 8'd21};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd244, 8'd158, 8'd49};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd241, 8'd171, 8'd39};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd251, 8'd181, 8'd51};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd254, 8'd166, 8'd66};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd212, 8'd107, 8'd41};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd37};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd188, 8'd80, 8'd44};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd182, 8'd102, 8'd43};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd160, 8'd57, 8'd22};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd142, 8'd24, 8'd0};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd157, 8'd51, 8'd0};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd154, 8'd81, 8'd28};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd190, 8'd152, 8'd141};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd192, 8'd185, 8'd193};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd167, 8'd179, 8'd179};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd178, 8'd186, 8'd188};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd180, 8'd204, 8'd206};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd161, 8'd189, 8'd190};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd145, 8'd144, 8'd139};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd121, 8'd73, 8'd53};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd131, 8'd40, 8'd9};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd177, 8'd71, 8'd31};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd159, 8'd56, 8'd15};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd147, 8'd47, 8'd0};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd176, 8'd79, 8'd34};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd174, 8'd77, 8'd35};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd161, 8'd55, 8'd13};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd186, 8'd74, 8'd28};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd203, 8'd91, 8'd51};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd155, 8'd57, 8'd32};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd90, 8'd7, 8'd0};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd136, 8'd51, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd203, 8'd105, 8'd70};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd179, 8'd64, 8'd19};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd178, 8'd60, 8'd12};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd191, 8'd80, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd175, 8'd71, 8'd32};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd166, 8'd60, 8'd20};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd183, 8'd72, 8'd29};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd195, 8'd78, 8'd34};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd189, 8'd77, 8'd37};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd168, 8'd61, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd149, 8'd49, 8'd17};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd143, 8'd43, 8'd11};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd195, 8'd88, 8'd52};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd192, 8'd80, 8'd40};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd188, 8'd71, 8'd27};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd176, 8'd71, 8'd26};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd164, 8'd55, 8'd12};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd171, 8'd58, 8'd16};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd185, 8'd69, 8'd28};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd185, 8'd69, 8'd28};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd184, 8'd71, 8'd29};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd185, 8'd76, 8'd33};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd179, 8'd74, 8'd29};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd155, 8'd44, 8'd0};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd179, 8'd71, 8'd25};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd160, 8'd61, 8'd22};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd120, 8'd36, 8'd10};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd96, 8'd30, 8'd16};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd112, 8'd50, 8'd37};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd146, 8'd71, 8'd48};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd144, 8'd58, 8'd23};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd144, 8'd52, 8'd31};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd141, 8'd57, 8'd29};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd121, 8'd43, 8'd7};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd128, 8'd46, 8'd9};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd133, 8'd42, 8'd11};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd131, 8'd41, 8'd17};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd96, 8'd19, 8'd1};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd85, 8'd19, 8'd3};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd130, 8'd50, 8'd23};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd152, 8'd69, 8'd39};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd138, 8'd52, 8'd19};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd142, 8'd50, 8'd13};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd132, 8'd38, 8'd0};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd142, 8'd48, 8'd10};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd141, 8'd49, 8'd12};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd127, 8'd35, 8'd0};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd155, 8'd102, 8'd70};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd192, 8'd187, 8'd184};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd158, 8'd187, 8'd203};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd127, 8'd154, 8'd163};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd114, 8'd135, 8'd140};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd122, 8'd146, 8'd158};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd146, 8'd156, 8'd165};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd168, 8'd151, 8'd144};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd147, 8'd62, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd174, 8'd86, 8'd23};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd188, 8'd98, 8'd36};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd178, 8'd88, 8'd28};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd159, 8'd66, 8'd9};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd145, 8'd49, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd152, 8'd54, 8'd5};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd171, 8'd73, 8'd26};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd235, 8'd161, 8'd26};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd251, 8'd183, 8'd48};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd241, 8'd171, 8'd47};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd83};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd230, 8'd100, 8'd51};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd213, 8'd50, 8'd33};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd220, 8'd42, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd215, 8'd50, 8'd46};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd222, 8'd54, 8'd51};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd230, 8'd61, 8'd58};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd237, 8'd63, 8'd62};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd237, 8'd57, 8'd58};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd230, 8'd46, 8'd48};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd219, 8'd33, 8'd36};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd213, 8'd24, 8'd28};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd208, 8'd23, 8'd20};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd211, 8'd16, 8'd12};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd206, 8'd19, 8'd12};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd193, 8'd20, 8'd13};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd201, 8'd17, 8'd17};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd205, 8'd12, 8'd5};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd211, 8'd63, 8'd17};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd82};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd245, 8'd175, 8'd43};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd32};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd249, 8'd185, 8'd79};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd192, 8'd123, 8'd84};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd214, 8'd149, 8'd107};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd221, 8'd159, 8'd110};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd104: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd240, 8'd204, 8'd180};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd234, 8'd187, 8'd159};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd227, 8'd176, 8'd147};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd192, 8'd141, 8'd112};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd183, 8'd133, 8'd106};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd171, 8'd95, 8'd61};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd216, 8'd125, 8'd54};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd45};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd146, 8'd21};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd63};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd224, 8'd97, 8'd44};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd188, 8'd21, 8'd3};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd236, 8'd33, 8'd36};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd204, 8'd19, 8'd24};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd203, 8'd20, 8'd24};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd206, 8'd23, 8'd27};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd215, 8'd35, 8'd38};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd230, 8'd50, 8'd53};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd238, 8'd59, 8'd62};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd240, 8'd61, 8'd64};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd238, 8'd59, 8'd62};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd226, 8'd66, 8'd66};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd222, 8'd57, 8'd51};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd229, 8'd55, 8'd46};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd222, 8'd38, 8'd38};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd234, 8'd48, 8'd59};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd219, 8'd39, 8'd48};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd212, 8'd43, 8'd38};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd193, 8'd32, 8'd12};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd243, 8'd154, 8'd70};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd250, 8'd167, 8'd47};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd234, 8'd159, 8'd6};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd242, 8'd165, 8'd27};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd245, 8'd160, 8'd70};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd159, 8'd67, 8'd16};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd145, 8'd52, 8'd8};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd179, 8'd88, 8'd33};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd167, 8'd87, 8'd18};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd175, 8'd70, 8'd12};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd189, 8'd61, 8'd14};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd182, 8'd56, 8'd16};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd180, 8'd87, 8'd53};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd201, 8'd154, 8'd128};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd197, 8'd190, 8'd174};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd171, 8'd184, 8'd175};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd166, 8'd179, 8'd185};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd177, 8'd188, 8'd194};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd170, 8'd196, 8'd195};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd123, 8'd153, 8'd141};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd128, 8'd110, 8'd96};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd138, 8'd51, 8'd34};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd171, 8'd61, 8'd28};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd161, 8'd72, 8'd16};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd156, 8'd49, 8'd17};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd186, 8'd78, 8'd40};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd169, 8'd58, 8'd13};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd161, 8'd51, 8'd2};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd174, 8'd67, 8'd21};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd187, 8'd88, 8'd47};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd176, 8'd85, 8'd54};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd112, 8'd26, 8'd1};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd135, 8'd44, 8'd23};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd198, 8'd100, 8'd71};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd189, 8'd82, 8'd40};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd185, 8'd71, 8'd19};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd193, 8'd76, 8'd23};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd189, 8'd74, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd167, 8'd59, 8'd21};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd170, 8'd67, 8'd36};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd200, 8'd79, 8'd36};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd185, 8'd72, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd172, 8'd72, 8'd36};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd145, 8'd55, 8'd21};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd131, 8'd40, 8'd9};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd173, 8'd73, 8'd41};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd211, 8'd97, 8'd61};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd197, 8'd75, 8'd38};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd184, 8'd81, 8'd38};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd171, 8'd65, 8'd23};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd169, 8'd60, 8'd19};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd192, 8'd79, 8'd39};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd186, 8'd73, 8'd33};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd188, 8'd79, 8'd38};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd177, 8'd71, 8'd29};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd168, 8'd65, 8'd22};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd11};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd10};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd149, 8'd65, 8'd29};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd111, 8'd35, 8'd11};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd84, 8'd9, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd119, 8'd41, 8'd19};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd147, 8'd60, 8'd33};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd142, 8'd47, 8'd17};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd137, 8'd45, 8'd20};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd144, 8'd61, 8'd31};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd137, 8'd61, 8'd27};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd131, 8'd51, 8'd18};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd133, 8'd43, 8'd17};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd120, 8'd29, 8'd8};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd95, 8'd18, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd84, 8'd22, 8'd1};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd124, 8'd47, 8'd37};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd151, 8'd61, 8'd27};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd130, 8'd42, 8'd2};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd137, 8'd62, 8'd33};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd122, 8'd35, 8'd8};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd149, 8'd40, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd143, 8'd46, 8'd4};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd112, 8'd48, 8'd21};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd145, 8'd129, 8'd114};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd186, 8'd182, 8'd170};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd166, 8'd183, 8'd177};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd123, 8'd162, 8'd169};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd117, 8'd163, 8'd176};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd119, 8'd144, 8'd151};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd164, 8'd150, 8'd139};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd173, 8'd127, 8'd101};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd173, 8'd66, 8'd34};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd191, 8'd85, 8'd46};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd191, 8'd86, 8'd38};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd165, 8'd60, 8'd3};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd147, 8'd40, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd153, 8'd45, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd167, 8'd55, 8'd18};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd169, 8'd56, 8'd26};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd220, 8'd130, 8'd34};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd38};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd245, 8'd164, 8'd21};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd243, 8'd187, 8'd48};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd246, 8'd157, 8'd67};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd211, 8'd45, 8'd19};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd237, 8'd42, 8'd40};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd225, 8'd48, 8'd42};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd223, 8'd54, 8'd49};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd227, 8'd55, 8'd51};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd230, 8'd55, 8'd52};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd230, 8'd50, 8'd49};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd226, 8'd40, 8'd41};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd216, 8'd26, 8'd28};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd206, 8'd11, 8'd15};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd199, 8'd3, 8'd7};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd217, 8'd19, 8'd16};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd198, 8'd10, 8'd1};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd196, 8'd12, 8'd4};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd193, 8'd7, 8'd12};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd205, 8'd18, 8'd29};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd207, 8'd34, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd208, 8'd64, 8'd27};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd252, 8'd135, 8'd68};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd246, 8'd173, 8'd34};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd247, 8'd159, 8'd25};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd50};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd214, 8'd134, 8'd61};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd251, 8'd204, 8'd176};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd105: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd246, 8'd217, 8'd213};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd241, 8'd202, 8'd197};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd236, 8'd193, 8'd187};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd211, 8'd167, 8'd164};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd207, 8'd166, 8'd164};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd194, 8'd116, 8'd78};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd210, 8'd123, 8'd46};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd251, 8'd151, 8'd37};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd148, 8'd24};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd57};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd212, 8'd85, 8'd34};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd201, 8'd35, 8'd19};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd225, 8'd29, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd194, 8'd10, 8'd12};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd197, 8'd13, 8'd15};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd200, 8'd16, 8'd18};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd202, 8'd18, 8'd20};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd204, 8'd21, 8'd23};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd215, 8'd32, 8'd34};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd232, 8'd49, 8'd51};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd245, 8'd62, 8'd64};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd227, 8'd61, 8'd61};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd227, 8'd56, 8'd49};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd233, 8'd54, 8'd47};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd227, 8'd41, 8'd42};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd233, 8'd47, 8'd58};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd219, 8'd44, 8'd49};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd205, 8'd45, 8'd31};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd205, 8'd56, 8'd24};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd252, 8'd168, 8'd70};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd41};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd242, 8'd163, 8'd18};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd242, 8'd160, 8'd34};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd201, 8'd110, 8'd31};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd147, 8'd50, 8'd5};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd138, 8'd40, 8'd0};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd156, 8'd60, 8'd2};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd171, 8'd88, 8'd48};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd201, 8'd100, 8'd56};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd190, 8'd73, 8'd20};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd166, 8'd54, 8'd0};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd182, 8'd101, 8'd36};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd195, 8'd157, 8'd108};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd182, 8'd181, 8'd160};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd179, 8'd199, 8'd198};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd172, 8'd185, 8'd191};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd183, 8'd192, 8'd199};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd184, 8'd204, 8'd205};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd132, 8'd158, 8'd149};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd131, 8'd113, 8'd101};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd134, 8'd48, 8'd33};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd166, 8'd57, 8'd26};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd159, 8'd68, 8'd15};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd152, 8'd48, 8'd13};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd181, 8'd75, 8'd35};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd164, 8'd56, 8'd10};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd159, 8'd51, 8'd2};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd173, 8'd67, 8'd19};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd187, 8'd85, 8'd45};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd182, 8'd85, 8'd53};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd123, 8'd31, 8'd6};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd131, 8'd39, 8'd16};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd197, 8'd98, 8'd67};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd188, 8'd81, 8'd39};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd182, 8'd66, 8'd15};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd188, 8'd71, 8'd17};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd189, 8'd74, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd169, 8'd60, 8'd21};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd166, 8'd61, 8'd29};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd197, 8'd74, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd183, 8'd70, 8'd28};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd171, 8'd69, 8'd31};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd144, 8'd51, 8'd17};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd131, 8'd38, 8'd5};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd173, 8'd70, 8'd37};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd207, 8'd93, 8'd57};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd195, 8'd71, 8'd33};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd183, 8'd77, 8'd35};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd169, 8'd62, 8'd20};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd168, 8'd56, 8'd16};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd191, 8'd75, 8'd36};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd185, 8'd69, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd188, 8'd76, 8'd36};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd176, 8'd69, 8'd27};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd167, 8'd61, 8'd19};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd169, 8'd63, 8'd13};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd154, 8'd55, 8'd13};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd149, 8'd63, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd111, 8'd33, 8'd10};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd86, 8'd11, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd123, 8'd42, 8'd21};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd150, 8'd60, 8'd34};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd143, 8'd48, 8'd18};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd133, 8'd41, 8'd16};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd139, 8'd55, 8'd27};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd136, 8'd60, 8'd28};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd137, 8'd56, 8'd26};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd138, 8'd48, 8'd22};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd117, 8'd29, 8'd9};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd95, 8'd18, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd89, 8'd27, 8'd6};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd129, 8'd51, 8'd39};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd156, 8'd63, 8'd29};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd134, 8'd45, 8'd3};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd139, 8'd62, 8'd32};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd125, 8'd35, 8'd8};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd149, 8'd40, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd141, 8'd45, 8'd3};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd114, 8'd53, 8'd25};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd164, 8'd150, 8'd137};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd186, 8'd182, 8'd171};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd153, 8'd169, 8'd166};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd116, 8'd154, 8'd163};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd120, 8'd163, 8'd179};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd124, 8'd148, 8'd158};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd170, 8'd156, 8'd147};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd178, 8'd132, 8'd108};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd196, 8'd98, 8'd53};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd176, 8'd77, 8'd35};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd159, 8'd58, 8'd16};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd153, 8'd52, 8'd8};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd153, 8'd51, 8'd2};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd151, 8'd50, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd157, 8'd57, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd168, 8'd66, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd193, 8'd101, 8'd16};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd240, 8'd138, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd238, 8'd155, 8'd17};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd232, 8'd174, 8'd31};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd243, 8'd155, 8'd57};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd215, 8'd59, 8'd19};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd210, 8'd21, 8'd15};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd220, 8'd42, 8'd40};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd212, 8'd34, 8'd32};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd210, 8'd32, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd207, 8'd27, 8'd26};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd206, 8'd22, 8'd22};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd205, 8'd17, 8'd18};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd204, 8'd14, 8'd16};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd206, 8'd13, 8'd16};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd207, 8'd12, 8'd16};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd204, 8'd9, 8'd5};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd194, 8'd6, 8'd0};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd198, 8'd15, 8'd9};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd203, 8'd17, 8'd20};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd215, 8'd28, 8'd39};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd214, 8'd40, 8'd39};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd211, 8'd64, 8'd31};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd246, 8'd123, 8'd63};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd242, 8'd164, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd243, 8'd155, 8'd22};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd244, 8'd148, 8'd35};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd197, 8'd119, 8'd44};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd238, 8'd191, 8'd163};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd106: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd213, 8'd132, 8'd85};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd206, 8'd120, 8'd37};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd237, 8'd144, 8'd25};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd248, 8'd150, 8'd27};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd253, 8'd145, 8'd55};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd197, 8'd66, 8'd20};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd213, 8'd50, 8'd35};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd220, 8'd32, 8'd31};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd193, 8'd8, 8'd6};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd194, 8'd9, 8'd7};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd193, 8'd8, 8'd6};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd191, 8'd6, 8'd4};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd192, 8'd7, 8'd5};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd203, 8'd18, 8'd16};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd220, 8'd35, 8'd33};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd233, 8'd48, 8'd46};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd225, 8'd51, 8'd50};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd44};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd235, 8'd47, 8'd45};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd232, 8'd41, 8'd46};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd226, 8'd41, 8'd49};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd216, 8'd48, 8'd45};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd194, 8'd46, 8'd18};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd225, 8'd91, 8'd40};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd255, 8'd178, 8'd60};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd245, 8'd164, 8'd31};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd247, 8'd165, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd234, 8'd146, 8'd38};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd161, 8'd64, 8'd0};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd149, 8'd46, 8'd5};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd146, 8'd41, 8'd0};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd149, 8'd45, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd156, 8'd66, 8'd40};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd174, 8'd76, 8'd39};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd196, 8'd91, 8'd33};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd185, 8'd89, 8'd5};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd167, 8'd96, 8'd6};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd189, 8'd154, 8'd88};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd209, 8'd208, 8'd187};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd185, 8'd204, 8'd218};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd182, 8'd195, 8'd201};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd195, 8'd197, 8'd209};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd222};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd146, 8'd167, 8'd162};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd137, 8'd120, 8'd110};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd127, 8'd48, 8'd33};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd158, 8'd50, 8'd21};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd158, 8'd63, 8'd15};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd147, 8'd48, 8'd7};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd175, 8'd74, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd160, 8'd55, 8'd7};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd160, 8'd54, 8'd4};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd174, 8'd68, 8'd20};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd187, 8'd81, 8'd41};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd189, 8'd86, 8'd55};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd144, 8'd42, 8'd17};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd129, 8'd33, 8'd8};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd197, 8'd97, 8'd65};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd190, 8'd81, 8'd38};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd178, 8'd62, 8'd11};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd182, 8'd65, 8'd12};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd192, 8'd76, 8'd27};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd175, 8'd63, 8'd23};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd164, 8'd56, 8'd20};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd193, 8'd71, 8'd24};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd183, 8'd68, 8'd24};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd170, 8'd66, 8'd27};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd145, 8'd48, 8'd13};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd134, 8'd37, 8'd4};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd172, 8'd68, 8'd33};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd205, 8'd89, 8'd52};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd193, 8'd70, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd182, 8'd75, 8'd31};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd168, 8'd59, 8'd16};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd167, 8'd54, 8'd12};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd189, 8'd73, 8'd32};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd183, 8'd67, 8'd26};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd186, 8'd73, 8'd31};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd174, 8'd65, 8'd22};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd166, 8'd59, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd170, 8'd62, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd157, 8'd55, 8'd15};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd149, 8'd60, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd111, 8'd30, 8'd9};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd90, 8'd13, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd128, 8'd46, 8'd25};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd34};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd147, 8'd49, 8'd20};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd128, 8'd38, 8'd14};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd129, 8'd48, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd130, 8'd55, 8'd23};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd142, 8'd61, 8'd31};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd145, 8'd58, 8'd31};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd120, 8'd32, 8'd12};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd94, 8'd19, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd92, 8'd31, 8'd12};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd138, 8'd56, 8'd45};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd163, 8'd66, 8'd31};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd141, 8'd48, 8'd4};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd143, 8'd63, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd128, 8'd37, 8'd6};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd149, 8'd40, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd137, 8'd44, 8'd1};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd118, 8'd62, 8'd35};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd171, 8'd161, 8'd151};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd192, 8'd189, 8'd182};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd157, 8'd173, 8'd173};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd113, 8'd149, 8'd161};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd114, 8'd155, 8'd175};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd121, 8'd143, 8'd156};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd166, 8'd151, 8'd144};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd165, 8'd119, 8'd96};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd169, 8'd83, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd181, 8'd91, 8'd13};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd181, 8'd89, 8'd24};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd170, 8'd75, 8'd19};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd164, 8'd67, 8'd14};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd169, 8'd73, 8'd13};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd173, 8'd76, 8'd8};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd168, 8'd72, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd176, 8'd79, 8'd8};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd221, 8'd119, 8'd21};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd235, 8'd148, 8'd15};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd230, 8'd164, 8'd18};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd41};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd228, 8'd89, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd183, 8'd10, 8'd0};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd208, 8'd32, 8'd34};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd203, 8'd15, 8'd16};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd200, 8'd12, 8'd13};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd196, 8'd6, 8'd8};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd192, 8'd2, 8'd4};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd192, 8'd2, 8'd4};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd195, 8'd5, 8'd7};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd199, 8'd9, 8'd11};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd202, 8'd12, 8'd14};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd198, 8'd3, 8'd1};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd193, 8'd6, 8'd0};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd203, 8'd22, 8'd15};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd213, 8'd30, 8'd32};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd224, 8'd38, 8'd49};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd46};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd212, 8'd61, 8'd34};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd234, 8'd105, 8'd50};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd249, 8'd163, 8'd40};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd250, 8'd158, 8'd31};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd240, 8'd146, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd196, 8'd119, 8'd39};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd227, 8'd178, 8'd146};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd107: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd210, 8'd124, 8'd67};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd209, 8'd124, 8'd33};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd227, 8'd141, 8'd18};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd248, 8'd153, 8'd33};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd143, 8'd61};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd187, 8'd49, 8'd12};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd216, 8'd52, 8'd42};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd225, 8'd46, 8'd42};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd207, 8'd20, 8'd15};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd200, 8'd13, 8'd8};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd194, 8'd7, 8'd2};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd195, 8'd6, 8'd2};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd202, 8'd13, 8'd9};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd207, 8'd18, 8'd14};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd210, 8'd18, 8'd15};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd209, 8'd17, 8'd14};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd217, 8'd33, 8'd33};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd223, 8'd34, 8'd32};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd231, 8'd35, 8'd36};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd231, 8'd36, 8'd44};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd214, 8'd29, 8'd37};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd207, 8'd45, 8'd34};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd188, 8'd53, 8'd6};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd239, 8'd123, 8'd50};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd40};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd238, 8'd158, 8'd19};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd242, 8'd158, 8'd33};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd212, 8'd119, 8'd24};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd159, 8'd56, 8'd0};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd172, 8'd65, 8'd19};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd170, 8'd63, 8'd9};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd165, 8'd58, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd155, 8'd60, 8'd4};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd156, 8'd59, 8'd6};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd183, 8'd87, 8'd27};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd188, 8'd96, 8'd23};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd158, 8'd81, 8'd3};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd190, 8'd141, 8'd83};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd229, 8'd215, 8'd202};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd191, 8'd199, 8'd222};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd192, 8'd207, 8'd212};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd205, 8'd218};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd223, 8'd225, 8'd237};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd166, 8'd182, 8'd181};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd141, 8'd131, 8'd121};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd127, 8'd58, 8'd43};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd149, 8'd47, 8'd22};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd158, 8'd63, 8'd19};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd149, 8'd52, 8'd9};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd171, 8'd73, 8'd26};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd158, 8'd58, 8'd9};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd162, 8'd60, 8'd11};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd175, 8'd70, 8'd25};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd185, 8'd79, 8'd40};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd197, 8'd90, 8'd58};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd166, 8'd58, 8'd32};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd129, 8'd31, 8'd4};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd198, 8'd95, 8'd62};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd192, 8'd85, 8'd43};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd175, 8'd63, 8'd13};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd178, 8'd62, 8'd11};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd195, 8'd80, 8'd33};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd183, 8'd70, 8'd28};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd164, 8'd54, 8'd17};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd187, 8'd69, 8'd21};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd183, 8'd70, 8'd26};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd173, 8'd67, 8'd28};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd147, 8'd47, 8'd13};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd140, 8'd40, 8'd8};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd176, 8'd69, 8'd35};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd201, 8'd87, 8'd50};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd190, 8'd71, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd182, 8'd75, 8'd31};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd168, 8'd59, 8'd16};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd167, 8'd54, 8'd12};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd190, 8'd72, 8'd32};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd184, 8'd66, 8'd26};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd187, 8'd74, 8'd32};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd175, 8'd66, 8'd23};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd167, 8'd60, 8'd16};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd168, 8'd59, 8'd18};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd157, 8'd54, 8'd21};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd145, 8'd55, 8'd29};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd108, 8'd27, 8'd10};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd16, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd131, 8'd48, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd151, 8'd59, 8'd34};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd147, 8'd49, 8'd20};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd39, 8'd15};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd119, 8'd38, 8'd11};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd118, 8'd43, 8'd12};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd140, 8'd61, 8'd31};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd154, 8'd66, 8'd42};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd127, 8'd40, 8'd21};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd94, 8'd18, 8'd2};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd88, 8'd27, 8'd8};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd142, 8'd60, 8'd49};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd165, 8'd68, 8'd33};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd146, 8'd50, 8'd2};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd144, 8'd62, 8'd25};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd129, 8'd39, 8'd5};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd147, 8'd42, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd129, 8'd44, 8'd3};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd124, 8'd77, 8'd51};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd178, 8'd171, 8'd165};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd195, 8'd196, 8'd191};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd159, 8'd174, 8'd179};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd113, 8'd146, 8'd161};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd112, 8'd150, 8'd171};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd124, 8'd144, 8'd155};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd161, 8'd144, 8'd136};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd139, 8'd93, 8'd67};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd179, 8'd99, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd204, 8'd122, 8'd10};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd211, 8'd126, 8'd19};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd189, 8'd101, 8'd3};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd179, 8'd85, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd195, 8'd95, 8'd20};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd209, 8'd105, 8'd42};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd208, 8'd102, 8'd44};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd188, 8'd89, 8'd21};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd205, 8'd104, 8'd12};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd236, 8'd144, 8'd17};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd241, 8'd162, 8'd17};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd28};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd246, 8'd127, 8'd45};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd179, 8'd24, 8'd0};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd190, 8'd14, 8'd16};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd203, 8'd4, 8'd9};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd203, 8'd4, 8'd9};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd200, 8'd4, 8'd8};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd198, 8'd3, 8'd7};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd194, 8'd4, 8'd6};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd193, 8'd5, 8'd6};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd191, 8'd5, 8'd6};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd191, 8'd5, 8'd6};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd207, 8'd13, 8'd14};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd200, 8'd17, 8'd11};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd207, 8'd30, 8'd22};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd217, 8'd39, 8'd39};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd226, 8'd40, 8'd51};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd220, 8'd41, 8'd45};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd213, 8'd56, 8'd37};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd221, 8'd84, 8'd40};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd56};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd250, 8'd153, 8'd36};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd240, 8'd150, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd207, 8'd130, 8'd40};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd207, 8'd152, 8'd111};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd108: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd198, 8'd101, 8'd33};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd221, 8'd133, 8'd35};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd229, 8'd145, 8'd20};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd250, 8'd155, 8'd39};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd255, 8'd139, 8'd68};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd185, 8'd37, 8'd11};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd211, 8'd44, 8'd38};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd235, 8'd62, 8'd58};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd216, 8'd33, 8'd27};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd209, 8'd24, 8'd19};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd200, 8'd15, 8'd10};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd198, 8'd11, 8'd6};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd199, 8'd10, 8'd6};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd201, 8'd9, 8'd6};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd197, 8'd3, 8'd1};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd192, 8'd0, 8'd0};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd204, 8'd16, 8'd14};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd212, 8'd18, 8'd16};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd220, 8'd20, 8'd23};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd224, 8'd23, 8'd33};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd201, 8'd14, 8'd21};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd195, 8'd39, 8'd17};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd192, 8'd68, 8'd4};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd246, 8'd144, 8'd46};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd249, 8'd169, 8'd22};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd234, 8'd152, 8'd14};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd230, 8'd144, 8'd25};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd186, 8'd93, 8'd0};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd180, 8'd81, 8'd13};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd193, 8'd91, 8'd29};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd187, 8'd84, 8'd17};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd182, 8'd79, 8'd2};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd179, 8'd84, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd189, 8'd98, 8'd19};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd169, 8'd82, 8'd29};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd164, 8'd73, 8'd28};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd168, 8'd80, 8'd34};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd184, 8'd116, 8'd81};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd210, 8'd176, 8'd174};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd203, 8'd197, 8'd223};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd194, 8'd213, 8'd217};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd211, 8'd207, 8'd221};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd228, 8'd226, 8'd239};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd180, 8'd196, 8'd196};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd141, 8'd141, 8'd131};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd130, 8'd74, 8'd59};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd136, 8'd44, 8'd19};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd155, 8'd63, 8'd24};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd151, 8'd56, 8'd10};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd169, 8'd74, 8'd28};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd155, 8'd60, 8'd14};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd162, 8'd67, 8'd21};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd170, 8'd73, 8'd31};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd174, 8'd74, 8'd38};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd194, 8'd91, 8'd60};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd179, 8'd74, 8'd45};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd131, 8'd32, 8'd3};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd194, 8'd94, 8'd62};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd189, 8'd85, 8'd46};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd174, 8'd67, 8'd21};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd173, 8'd62, 8'd16};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd194, 8'd83, 8'd38};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd187, 8'd75, 8'd35};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd168, 8'd56, 8'd19};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd181, 8'd69, 8'd21};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd183, 8'd74, 8'd31};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd172, 8'd68, 8'd31};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd148, 8'd47, 8'd17};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd144, 8'd43, 8'd13};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd176, 8'd71, 8'd39};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd196, 8'd86, 8'd49};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd186, 8'd73, 8'd33};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd182, 8'd76, 8'd34};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd168, 8'd61, 8'd19};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd167, 8'd55, 8'd15};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd188, 8'd75, 8'd35};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd182, 8'd69, 8'd29};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd187, 8'd75, 8'd35};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd175, 8'd68, 8'd26};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd167, 8'd61, 8'd19};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd164, 8'd56, 8'd18};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd151, 8'd52, 8'd21};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd137, 8'd49, 8'd27};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd99, 8'd22, 8'd6};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd17, 8'd4};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd131, 8'd50, 8'd33};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd145, 8'd57, 8'd33};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd144, 8'd49, 8'd19};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd129, 8'd41, 8'd19};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd112, 8'd32, 8'd5};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd104, 8'd31, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd130, 8'd53, 8'd23};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd155, 8'd69, 8'd46};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd133, 8'd46, 8'd27};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd93, 8'd20, 8'd3};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd78, 8'd19, 8'd1};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd140, 8'd60, 8'd51};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd162, 8'd65, 8'd32};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd144, 8'd49, 8'd3};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd141, 8'd59, 8'd22};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd127, 8'd38, 8'd4};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd144, 8'd43, 8'd0};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd122, 8'd44, 8'd6};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd129, 8'd93, 8'd71};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd190, 8'd188, 8'd189};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd185, 8'd189, 8'd192};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd147, 8'd161, 8'd170};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd116, 8'd147, 8'd165};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd119, 8'd154, 8'd173};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd128, 8'd145, 8'd152};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd172, 8'd157, 8'd138};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd161, 8'd119, 8'd81};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd234, 8'd158, 8'd83};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd219, 8'd144, 8'd53};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd210, 8'd133, 8'd19};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd214, 8'd133, 8'd2};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd220, 8'd132, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd221, 8'd125, 8'd5};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd224, 8'd117, 8'd19};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd227, 8'd117, 8'd32};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd217, 8'd118, 8'd37};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd196, 8'd99, 8'd2};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd232, 8'd138, 8'd16};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd251, 8'd160, 8'd19};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd235, 8'd152, 8'd14};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd249, 8'd153, 8'd50};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd191, 8'd56, 8'd8};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd171, 8'd0, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd202, 8'd1, 8'd7};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd202, 8'd1, 8'd7};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd199, 8'd3, 8'd7};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd199, 8'd4, 8'd8};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd198, 8'd8, 8'd10};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd199, 8'd11, 8'd12};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd198, 8'd14, 8'd14};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd199, 8'd15, 8'd15};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd226, 8'd33, 8'd36};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd216, 8'd34, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd211, 8'd39, 8'd29};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd219, 8'd35, 8'd45};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd215, 8'd34, 8'd43};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd214, 8'd50, 8'd40};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd211, 8'd64, 8'd31};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd255, 8'd144, 8'd64};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd246, 8'd141, 8'd36};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd236, 8'd144, 8'd21};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd214, 8'd133, 8'd28};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd184, 8'd118, 8'd60};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd248, 8'd206, 8'd192};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd109: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd244, 8'd209, 8'd205};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd200, 8'd92, 8'd17};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd234, 8'd141, 8'd37};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd233, 8'd150, 8'd22};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd253, 8'd155, 8'd44};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd251, 8'd121, 8'd59};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd191, 8'd31, 8'd15};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd207, 8'd35, 8'd35};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd239, 8'd67, 8'd65};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd218, 8'd39, 8'd35};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd216, 8'd37, 8'd33};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd211, 8'd29, 8'd26};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd200, 8'd15, 8'd13};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd189, 8'd1, 8'd0};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd184, 8'd0, 8'd0};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd190, 8'd0, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd196, 8'd2, 8'd3};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd193, 8'd6, 8'd0};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd202, 8'd7, 8'd3};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd211, 8'd6, 8'd11};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd216, 8'd12, 8'd24};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd193, 8'd4, 8'd10};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd188, 8'd33, 8'd5};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd214, 8'd94, 8'd16};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd248, 8'd154, 8'd38};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd244, 8'd159, 8'd14};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd234, 8'd147, 8'd14};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd218, 8'd129, 8'd13};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd180, 8'd91, 8'd0};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd204, 8'd113, 8'd22};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd200, 8'd108, 8'd21};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd193, 8'd101, 8'd14};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd190, 8'd98, 8'd11};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd181, 8'd98, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd196, 8'd124, 8'd40};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd196, 8'd129, 8'd86};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd199, 8'd124, 8'd93};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd175, 8'd91, 8'd55};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd165, 8'd92, 8'd59};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd204, 8'd163, 8'd157};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd212, 8'd200, 8'd222};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd182, 8'd210, 8'd211};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd202, 8'd200, 8'd214};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd217, 8'd210, 8'd226};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd185, 8'd203, 8'd205};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd132, 8'd142, 8'd131};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd131, 8'd92, 8'd75};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd120, 8'd40, 8'd15};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd146, 8'd61, 8'd24};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd152, 8'd55, 8'd13};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd163, 8'd70, 8'd27};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd148, 8'd56, 8'd15};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd156, 8'd68, 8'd28};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd157, 8'd69, 8'd31};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd154, 8'd64, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd181, 8'd86, 8'd56};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd179, 8'd81, 8'd54};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd127, 8'd31, 8'd6};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd183, 8'd85, 8'd56};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd180, 8'd82, 8'd47};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd171, 8'd69, 8'd29};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd166, 8'd63, 8'd22};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd185, 8'd79, 8'd39};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd182, 8'd74, 8'd36};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd166, 8'd58, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd172, 8'd65, 8'd21};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd177, 8'd73, 8'd34};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd166, 8'd66, 8'd34};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd142, 8'd44, 8'd17};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd143, 8'd45, 8'd20};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd171, 8'd70, 8'd42};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd186, 8'd81, 8'd49};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd179, 8'd71, 8'd33};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd174, 8'd75, 8'd36};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd161, 8'd59, 8'd21};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd160, 8'd53, 8'd17};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd182, 8'd72, 8'd37};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd176, 8'd66, 8'd31};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd180, 8'd73, 8'd37};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd168, 8'd66, 8'd28};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd159, 8'd60, 8'd21};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd154, 8'd51, 8'd18};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd145, 8'd50, 8'd22};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd126, 8'd44, 8'd23};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd88, 8'd14, 8'd1};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd88, 8'd18, 8'd6};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd126, 8'd51, 8'd32};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd139, 8'd55, 8'd29};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd137, 8'd48, 8'd16};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd126, 8'd39, 8'd19};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd109, 8'd32, 8'd6};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd100, 8'd26, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd120, 8'd43, 8'd15};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd146, 8'd60, 8'd37};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd130, 8'd44, 8'd27};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd90, 8'd18, 8'd3};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd72, 8'd13, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd133, 8'd55, 8'd51};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd153, 8'd60, 8'd29};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd138, 8'd45, 8'd1};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd134, 8'd54, 8'd19};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd122, 8'd38, 8'd4};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd138, 8'd45, 8'd4};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd112, 8'd46, 8'd12};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd132, 8'd109, 8'd95};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd184, 8'd184, 8'd194};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd170, 8'd174, 8'd185};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd141, 8'd157, 8'd170};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd126, 8'd155, 8'd171};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd115, 8'd147, 8'd160};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd116, 8'd133, 8'd127};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd198, 8'd184, 8'd149};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd236, 8'd197, 8'd140};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd194};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd248, 8'd190, 8'd152};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd225, 8'd163, 8'd86};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd213, 8'd146, 8'd31};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd220, 8'd145, 8'd2};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd233, 8'd148, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd236, 8'd142, 8'd0};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd231, 8'd131, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd238, 8'd142, 8'd32};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd201, 8'd110, 8'd0};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd229, 8'd130, 8'd10};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd251, 8'd148, 8'd17};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd231, 8'd145, 8'd6};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd237, 8'd163, 8'd42};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd211, 8'd96, 8'd29};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd169, 8'd0, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd201, 8'd5, 8'd9};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd199, 8'd4, 8'd8};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd198, 8'd3, 8'd7};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd197, 8'd7, 8'd9};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd202, 8'd14, 8'd15};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd209, 8'd23, 8'd24};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd216, 8'd32, 8'd32};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd221, 8'd39, 8'd38};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd238, 8'd47, 8'd54};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd226, 8'd49, 8'd43};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd213, 8'd45, 8'd34};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd216, 8'd44, 8'd40};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd213, 8'd31, 8'd43};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd211, 8'd29, 8'd41};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd217, 8'd48, 8'd43};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd204, 8'd48, 8'd26};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd248, 8'd119, 8'd64};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd144, 8'd52};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd242, 8'd144, 8'd19};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd228, 8'd137, 8'd20};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd192, 8'd109, 8'd33};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd236, 8'd173, 8'd140};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd110: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd241, 8'd242, 8'd224};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd210};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd255, 8'd223, 8'd185};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd206, 8'd157, 8'd116};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd228, 8'd109, 8'd27};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd242, 8'd144, 8'd35};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd237, 8'd152, 8'd25};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd50};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd230, 8'd90, 8'd37};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd201, 8'd30, 8'd22};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd212, 8'd33, 8'd37};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd231, 8'd59, 8'd59};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd217, 8'd43, 8'd42};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd218, 8'd40, 8'd40};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd212, 8'd29, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd200, 8'd16, 8'd18};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd195, 8'd6, 8'd10};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd196, 8'd5, 8'd10};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd200, 8'd7, 8'd12};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd186, 8'd2, 8'd0};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd196, 8'd3, 8'd0};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd205, 8'd0, 8'd7};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd211, 8'd4, 8'd20};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd191, 8'd0, 8'd7};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd187, 8'd30, 8'd0};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd241, 8'd126, 8'd37};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd249, 8'd161, 8'd28};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd241, 8'd151, 8'd15};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd232, 8'd143, 8'd15};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd211, 8'd122, 8'd4};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd208, 8'd123, 8'd7};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd222, 8'd138, 8'd24};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd211, 8'd131, 8'd18};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd208, 8'd129, 8'd26};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd209, 8'd130, 8'd35};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd193, 8'd128, 8'd46};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd203, 8'd156, 8'd100};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd230, 8'd194, 8'd160};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd253, 8'd208, 8'd166};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd197, 8'd136, 8'd73};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd158, 8'd98, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd201, 8'd166, 8'd144};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd200, 8'd196, 8'd211};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd164, 8'd200, 8'd198};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd186, 8'd185, 8'd199};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd194, 8'd187, 8'd203};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd182, 8'd201, 8'd205};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd117, 8'd137, 8'd125};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd130, 8'd104, 8'd87};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd101, 8'd31, 8'd6};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd136, 8'd53, 8'd19};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd148, 8'd50, 8'd13};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd155, 8'd61, 8'd25};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd136, 8'd51, 8'd14};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd143, 8'd63, 8'd28};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd140, 8'd61, 8'd28};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd131, 8'd50, 8'd20};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd161, 8'd78, 8'd48};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd168, 8'd81, 8'd54};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd120, 8'd28, 8'd5};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd168, 8'd74, 8'd48};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd166, 8'd73, 8'd42};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd163, 8'd69, 8'd35};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd156, 8'd60, 8'd22};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd171, 8'd71, 8'd35};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd171, 8'd68, 8'd33};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd159, 8'd54, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd156, 8'd57, 8'd16};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd167, 8'd69, 8'd34};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd155, 8'd60, 8'd32};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd133, 8'd37, 8'd15};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd136, 8'd39, 8'd20};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd160, 8'd64, 8'd40};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd173, 8'd74, 8'd43};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd166, 8'd66, 8'd32};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd163, 8'd69, 8'd33};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd150, 8'd53, 8'd18};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd148, 8'd48, 8'd14};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd171, 8'd66, 8'd34};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd165, 8'd60, 8'd28};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd168, 8'd68, 8'd34};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd156, 8'd59, 8'd24};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd147, 8'd53, 8'd17};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd145, 8'd48, 8'd16};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd137, 8'd47, 8'd21};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd115, 8'd38, 8'd20};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd78, 8'd10, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd84, 8'd18, 8'd4};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd120, 8'd52, 8'd33};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd129, 8'd52, 8'd24};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd131, 8'd47, 8'd13};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd118, 8'd31, 8'd11};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd113, 8'd36, 8'd10};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd104, 8'd33, 8'd5};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd112, 8'd37, 8'd8};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd130, 8'd45, 8'd24};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd117, 8'd34, 8'd16};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd87, 8'd15, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd71, 8'd14, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd122, 8'd50, 8'd51};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd143, 8'd53, 8'd26};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd130, 8'd41, 8'd0};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd125, 8'd49, 8'd15};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd116, 8'd37, 8'd6};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd131, 8'd46, 8'd9};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd104, 8'd47, 8'd18};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd134, 8'd121, 8'd112};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd163, 8'd166, 8'd183};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd155, 8'd161, 8'd177};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd133, 8'd149, 8'd164};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd115, 8'd143, 8'd157};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd103, 8'd134, 8'd139};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd118, 8'd135, 8'd117};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd219, 8'd207, 8'd157};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd154};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd214};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd212};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd250, 8'd217, 8'd172};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd214, 8'd169, 8'd102};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd205, 8'd146, 8'd52};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd229, 8'd160, 8'd33};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd252, 8'd172, 8'd21};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd251, 8'd168, 8'd0};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd248, 8'd155, 8'd15};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd227, 8'd140, 8'd7};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd231, 8'd131, 8'd11};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd250, 8'd137, 8'd15};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd239, 8'd153, 8'd18};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd227, 8'd167, 8'd35};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd237, 8'd137, 8'd52};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd199, 8'd30, 8'd0};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd208, 8'd20, 8'd21};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd210, 8'd22, 8'd23};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd210, 8'd24, 8'd25};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd214, 8'd28, 8'd29};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd220, 8'd34, 8'd35};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd226, 8'd42, 8'd42};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd232, 8'd48, 8'd48};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd235, 8'd51, 8'd51};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd239, 8'd50, 8'd57};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd227, 8'd52, 8'd47};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd212, 8'd48, 8'd36};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd218, 8'd51, 8'd45};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd215, 8'd35, 8'd46};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd215, 8'd30, 8'd44};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd223, 8'd49, 8'd51};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd200, 8'd36, 8'd24};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd215, 8'd72, 8'd38};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd74};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd251, 8'd147, 8'd22};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd243, 8'd142, 8'd12};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd223, 8'd123, 8'd29};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd215, 8'd134, 8'd79};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd171};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd214};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd111: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd226, 8'd228, 8'd163};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd237, 8'd220, 8'd142};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd232, 8'd192, 8'd104};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd162, 8'd108, 8'd12};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd254, 8'd129, 8'd45};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd246, 8'd144, 8'd33};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd238, 8'd153, 8'd24};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd155, 8'd52};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd211, 8'd65, 8'd16};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd207, 8'd29, 8'd25};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd217, 8'd36, 8'd43};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd220, 8'd48, 8'd48};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd218, 8'd48, 8'd48};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd219, 8'd47, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd220, 8'd46, 8'd47};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd225, 8'd46, 8'd49};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd228, 8'd45, 8'd49};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd221, 8'd35, 8'd40};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd207, 8'd18, 8'd24};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd196, 8'd5, 8'd12};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd184, 8'd4, 8'd0};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd195, 8'd3, 8'd0};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd204, 8'd0, 8'd6};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd210, 8'd2, 8'd18};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd192, 8'd1, 8'd8};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd187, 8'd30, 8'd0};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd255, 8'd146, 8'd51};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd252, 8'd162, 8'd22};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd238, 8'd145, 8'd16};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd231, 8'd139, 8'd16};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd210, 8'd121, 8'd1};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd241, 8'd157, 8'd33};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd231, 8'd154, 8'd22};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd222, 8'd152, 8'd22};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd229, 8'd159, 8'd45};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd231, 8'd162, 8'd61};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd232, 8'd180, 8'd143};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd250, 8'd220, 8'd194};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd231, 8'd220, 8'd190};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd249, 8'd231, 8'd169};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd236, 8'd196, 8'd101};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd172, 8'd126, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd167, 8'd145, 8'd106};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd183, 8'd187, 8'd198};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd150, 8'd190, 8'd189};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd170, 8'd174, 8'd186};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd176, 8'd169, 8'd187};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd175, 8'd199, 8'd201};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd105, 8'd131, 8'd118};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd127, 8'd110, 8'd92};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd86, 8'd24, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd125, 8'd46, 8'd13};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd145, 8'd45, 8'd11};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd149, 8'd55, 8'd21};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd128, 8'd44, 8'd10};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd134, 8'd58, 8'd26};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd127, 8'd53, 8'd24};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd114, 8'd40, 8'd11};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd146, 8'd69, 8'd41};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd158, 8'd78, 8'd51};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd115, 8'd24, 8'd3};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd155, 8'd65, 8'd41};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd154, 8'd64, 8'd37};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd156, 8'd67, 8'd35};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd149, 8'd56, 8'd23};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd161, 8'd64, 8'd31};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd162, 8'd62, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd155, 8'd52, 8'd21};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd145, 8'd52, 8'd11};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd159, 8'd65, 8'd31};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd148, 8'd54, 8'd29};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd124, 8'd31, 8'd13};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd128, 8'd35, 8'd18};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd153, 8'd58, 8'd38};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd162, 8'd67, 8'd39};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd155, 8'd60, 8'd28};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd153, 8'd63, 8'd29};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd142, 8'd47, 8'd15};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd140, 8'd43, 8'd11};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd162, 8'd61, 8'd31};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd155, 8'd54, 8'd24};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd159, 8'd62, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd148, 8'd53, 8'd21};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd138, 8'd48, 8'd14};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd140, 8'd45, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd131, 8'd45, 8'd20};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd108, 8'd35, 8'd18};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd71, 8'd7, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd80, 8'd18, 8'd5};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd117, 8'd52, 8'd32};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd124, 8'd50, 8'd21};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd126, 8'd46, 8'd11};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd111, 8'd24, 8'd5};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd117, 8'd39, 8'd16};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd111, 8'd40, 8'd12};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd109, 8'd33, 8'd7};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd117, 8'd32, 8'd11};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd106, 8'd23, 8'd7};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd85, 8'd13, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd73, 8'd16, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd115, 8'd46, 8'd49};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd135, 8'd49, 8'd24};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd126, 8'd38, 8'd0};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd120, 8'd47, 8'd15};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd112, 8'd37, 8'd8};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd127, 8'd47, 8'd12};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd100, 8'd49, 8'd22};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd134, 8'd129, 8'd123};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd154, 8'd159, 8'd179};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd146, 8'd153, 8'd172};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd113, 8'd129, 8'd145};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd87, 8'd113, 8'd126};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd98, 8'd129, 8'd131};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd144, 8'd162, 8'd136};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd230, 8'd220, 8'd158};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd232, 8'd198, 8'd111};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd204, 8'd228, 8'd142};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd234, 8'd246, 8'd180};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd178};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd243, 8'd181, 8'd108};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd235, 8'd165, 8'd51};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd237, 8'd165, 8'd21};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd252, 8'd163, 8'd1};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd254, 8'd169, 8'd26};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd241, 8'd138, 8'd17};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd250, 8'd133, 8'd19};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd253, 8'd166, 8'd33};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd223, 8'd171, 8'd35};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd69};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd232, 8'd65, 8'd23};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd219, 8'd37, 8'd36};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd225, 8'd43, 8'd42};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd234, 8'd52, 8'd51};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd241, 8'd59, 8'd58};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd245, 8'd61, 8'd61};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd242, 8'd58, 8'd58};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd237, 8'd53, 8'd53};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd233, 8'd49, 8'd49};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd233, 8'd43, 8'd53};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd225, 8'd50, 8'd45};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd213, 8'd49, 8'd37};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd223, 8'd56, 8'd50};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd220, 8'd40, 8'd51};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd219, 8'd34, 8'd50};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd227, 8'd50, 8'd56};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd197, 8'd30, 8'd21};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd171, 8'd20, 8'd1};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd79};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd249, 8'd141, 8'd15};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd243, 8'd137, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd242, 8'd131, 8'd26};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd187, 8'd94, 8'd27};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd199, 8'd149, 8'd98};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd223, 8'd211, 8'd159};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd112: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd239, 8'd217, 8'd157};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd202, 8'd137, 8'd53};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd199, 8'd99, 8'd5};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd228, 8'd122, 8'd10};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd243, 8'd136, 8'd20};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd37};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd255, 8'd127, 8'd62};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd180, 8'd33, 8'd15};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd192, 8'd28, 8'd37};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd216, 8'd43, 8'd47};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd41};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd212, 8'd31, 8'd20};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd202, 8'd19, 8'd11};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd211, 8'd26, 8'd24};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd202, 8'd22, 8'd25};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd184, 8'd22, 8'd11};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd215, 8'd85, 8'd33};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd247, 8'd152, 8'd42};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd230, 8'd159, 8'd9};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd20};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd242, 8'd149, 8'd10};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd232, 8'd146, 8'd11};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd228, 8'd152, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd226, 8'd162, 8'd62};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd228, 8'd179, 8'd103};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd246, 8'd208, 8'd159};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd202};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd255};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd253, 8'd223, 8'd215};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd232, 8'd216, 8'd156};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd230, 8'd216, 8'd109};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd242, 8'd217, 8'd101};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd240, 8'd208, 8'd125};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd220, 8'd185, 8'd163};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd197, 8'd167, 8'd191};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd167, 8'd166, 8'd161};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd161};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd155, 8'd154, 8'd168};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd171, 8'd180, 8'd195};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd120, 8'd131, 8'd135};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd116, 8'd109, 8'd99};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd81, 8'd43, 8'd20};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd94, 8'd29, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd106, 8'd48, 8'd28};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd125, 8'd59, 8'd33};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd110, 8'd37, 8'd5};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd139, 8'd69, 8'd43};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd122, 8'd61, 8'd43};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd88, 8'd30, 8'd18};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd130, 8'd65, 8'd47};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd146, 8'd71, 8'd48};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd122, 8'd46, 8'd23};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd106, 8'd30, 8'd6};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd137, 8'd59, 8'd36};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd136, 8'd59, 8'd33};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd135, 8'd55, 8'd28};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd137, 8'd56, 8'd29};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd140, 8'd59, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd129, 8'd45, 8'd17};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd127, 8'd50, 8'd22};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd132, 8'd56, 8'd32};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd127, 8'd55, 8'd31};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd97, 8'd29, 8'd8};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd104, 8'd36, 8'd15};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd142, 8'd70, 8'd46};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd144, 8'd68, 8'd44};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd134, 8'd57, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd138, 8'd57, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd129, 8'd48, 8'd21};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd124, 8'd44, 8'd17};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd130, 8'd50, 8'd23};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd131, 8'd54, 8'd26};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd125, 8'd50, 8'd21};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd121, 8'd46, 8'd17};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd122, 8'd47, 8'd18};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd103, 8'd35, 8'd12};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd105, 8'd43, 8'd22};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd97, 8'd40, 8'd21};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd64, 8'd13, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd69, 8'd18, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd106, 8'd49, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd108, 8'd46, 8'd25};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd99, 8'd31, 8'd8};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd91, 8'd27, 8'd15};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd85, 8'd29, 8'd12};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd83, 8'd33, 8'd10};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd90, 8'd33, 8'd13};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd98, 8'd33, 8'd15};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd94, 8'd28, 8'd14};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd76, 8'd22, 8'd10};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd60, 8'd18, 8'd4};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd85, 8'd40, 8'd19};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd114, 8'd58, 8'd35};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd107, 8'd37, 8'd11};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd111, 8'd36, 8'd7};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd104, 8'd37, 8'd11};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd83, 8'd38, 8'd17};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd71, 8'd53, 8'd39};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd141, 8'd141, 8'd131};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd157, 8'd135, 8'd181};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd133, 8'd132, 8'd138};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd97, 8'd118, 8'd113};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd81, 8'd109, 8'd130};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd80, 8'd102, 8'd123};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd157, 8'd166, 8'd137};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd254, 8'd242, 8'd166};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd236, 8'd210, 8'd115};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd242, 8'd217, 8'd54};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd242, 8'd220, 8'd109};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd247, 8'd230, 8'd186};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd207};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd247, 8'd211, 8'd159};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd234, 8'd188, 8'd129};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd239, 8'd173, 8'd63};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd243, 8'd155, 8'd49};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd248, 8'd140, 8'd31};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd239, 8'd135, 8'd10};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd237, 8'd154, 8'd14};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd239, 8'd162, 8'd34};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd255, 8'd160, 8'd68};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd220, 8'd104, 8'd45};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd219, 8'd60, 8'd38};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd249, 8'd56, 8'd57};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd252, 8'd52, 8'd65};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd227, 8'd57, 8'd58};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd220, 8'd62, 8'd51};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd234, 8'd55, 8'd48};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd239, 8'd48, 8'd53};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd232, 8'd52, 8'd61};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd227, 8'd51, 8'd51};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd215, 8'd39, 8'd39};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd213, 8'd37, 8'd37};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd193, 8'd20, 8'd13};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd215, 8'd80, 8'd32};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd62};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd224, 8'd135, 8'd5};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd234, 8'd134, 8'd12};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd212, 8'd116, 8'd29};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd188, 8'd128, 8'd76};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd204};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd113: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd249, 8'd218, 8'd171};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd193, 8'd115, 8'd41};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd221, 8'd106, 8'd17};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd229, 8'd128, 8'd12};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd245, 8'd140, 8'd23};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd255, 8'd143, 8'd44};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd227, 8'd94, 8'd35};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd183, 8'd31, 8'd17};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd201, 8'd34, 8'd44};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd217, 8'd40, 8'd48};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd228, 8'd49, 8'd42};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd235, 8'd54, 8'd47};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd229, 8'd45, 8'd43};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd234, 8'd50, 8'd52};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd224, 8'd45, 8'd48};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd211, 8'd54, 8'd35};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd243, 8'd117, 8'd58};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd255, 8'd173, 8'd62};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd242, 8'd170, 8'd23};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd229, 8'd150, 8'd23};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd227, 8'd155, 8'd37};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd228, 8'd169, 8'd69};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd240, 8'd194, 8'd116};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd168};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd248, 8'd240, 8'd157};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd231, 8'd228, 8'd133};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd221, 8'd221, 8'd107};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd233, 8'd228, 8'd98};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd254, 8'd239, 8'd110};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd252, 8'd234, 8'd132};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd219, 8'd210, 8'd151};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd184, 8'd187, 8'd160};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd155, 8'd152, 8'd161};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd144, 8'd137, 8'd155};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd146, 8'd141, 8'd171};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd157, 8'd160, 8'd191};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd117, 8'd122, 8'd142};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd110, 8'd100, 8'd108};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd88, 8'd49, 8'd44};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd102, 8'd38, 8'd26};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd98, 8'd39, 8'd9};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd116, 8'd48, 8'd13};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd105, 8'd30, 8'd0};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd127, 8'd54, 8'd19};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd115, 8'd54, 8'd26};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd78, 8'd20, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd122, 8'd56, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd135, 8'd60, 8'd28};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd117, 8'd41, 8'd9};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd101, 8'd25, 8'd0};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd132, 8'd53, 8'd20};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd130, 8'd51, 8'd18};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd127, 8'd47, 8'd12};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd131, 8'd49, 8'd12};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd134, 8'd52, 8'd15};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd121, 8'd39, 8'd1};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd120, 8'd42, 8'd4};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd123, 8'd47, 8'd13};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd120, 8'd47, 8'd15};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd92, 8'd21, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd98, 8'd27, 8'd0};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd134, 8'd61, 8'd29};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd135, 8'd59, 8'd25};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd126, 8'd48, 8'd10};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd131, 8'd49, 8'd12};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd121, 8'd39, 8'd2};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd116, 8'd36, 8'd0};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd121, 8'd41, 8'd4};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd123, 8'd45, 8'd7};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd116, 8'd41, 8'd2};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd112, 8'd37, 8'd0};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd114, 8'd39, 8'd0};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd100, 8'd26, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd100, 8'd32, 8'd23};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd92, 8'd32, 8'd24};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd62, 8'd5, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd67, 8'd10, 8'd3};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd100, 8'd40, 8'd32};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd104, 8'd36, 8'd27};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd96, 8'd22, 8'd11};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd88, 8'd23, 8'd1};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd81, 8'd24, 8'd0};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd78, 8'd28, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd85, 8'd29, 8'd0};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd94, 8'd27, 8'd0};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd90, 8'd22, 8'd0};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd72, 8'd17, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd55, 8'd13, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd81, 8'd35, 8'd2};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd115, 8'd56, 8'd22};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd110, 8'd40, 8'd4};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd110, 8'd34, 8'd0};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd102, 8'd33, 8'd0};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd77, 8'd30, 8'd4};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd82, 8'd61, 8'd42};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd134, 8'd131, 8'd116};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd123, 8'd133, 8'd145};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd96, 8'd121, 8'd102};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd80, 8'd119, 8'd98};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd79, 8'd117, 8'd126};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd88, 8'd115, 8'd124};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd165, 8'd174, 8'd131};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd254, 8'd241, 8'd149};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd119};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd251, 8'd217, 8'd128};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd239, 8'd216, 8'd122};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd227, 8'd220, 8'd130};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd234, 8'd235, 8'd175};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd241, 8'd240, 8'd194};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd245, 8'd221, 8'd147};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd249, 8'd200, 8'd131};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd248, 8'd177, 8'd99};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd230, 8'd155, 8'd54};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd226, 8'd156, 8'd34};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd230, 8'd156, 8'd35};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd66};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd245, 8'd124, 8'd53};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd219, 8'd65, 8'd39};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd246, 8'd57, 8'd55};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd250, 8'd52, 8'd65};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd228, 8'd58, 8'd61};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd220, 8'd62, 8'd51};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd234, 8'd55, 8'd48};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd240, 8'd49, 8'd54};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd231, 8'd51, 8'd60};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd227, 8'd51, 8'd51};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd215, 8'd39, 8'd39};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd213, 8'd37, 8'd37};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd201, 8'd27, 8'd20};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd202, 8'd61, 8'd18};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd251, 8'd146, 8'd55};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd232, 8'd136, 8'd15};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd235, 8'd131, 8'd10};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd223, 8'd126, 8'd32};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd185, 8'd120, 8'd64};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd244, 8'd211, 8'd178};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd114: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd237, 8'd194, 8'd160};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd197, 8'd102, 8'd34};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd246, 8'd112, 8'd23};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd232, 8'd136, 8'd15};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd252, 8'd148, 8'd35};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd247, 8'd129, 8'd41};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd191, 8'd55, 8'd5};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd186, 8'd29, 8'd20};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd210, 8'd38, 8'd50};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd218, 8'd36, 8'd48};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd229, 8'd45, 8'd47};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd241, 8'd59, 8'd58};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd242, 8'd57, 8'd62};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd243, 8'd60, 8'd65};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd230, 8'd57, 8'd53};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd228, 8'd77, 8'd48};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd68};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd63};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd233, 8'd165, 8'd22};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd210, 8'd158, 8'd57};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd237, 8'd196, 8'd114};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd180};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd233, 8'd217, 8'd95};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd235, 8'd218, 8'd102};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd243, 8'd219, 8'd109};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd113};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd113};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd247, 8'd208, 8'd115};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd214, 8'd197, 8'd125};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd186, 8'd189, 8'd132};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd142, 8'd145, 8'd150};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd118, 8'd116, 8'd130};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd123, 8'd121, 8'd145};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd129, 8'd133, 8'd160};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd114, 8'd121, 8'd140};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd101, 8'd96, 8'd102};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd79, 8'd48, 8'd43};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd78, 8'd26, 8'd15};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd92, 8'd32, 8'd22};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd104, 8'd37, 8'd21};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd102, 8'd27, 8'd6};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd111, 8'd39, 8'd24};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd111, 8'd48, 8'd41};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd72, 8'd12, 8'd11};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd118, 8'd51, 8'd43};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd124, 8'd50, 8'd37};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd113, 8'd39, 8'd26};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd97, 8'd21, 8'd8};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd125, 8'd49, 8'd35};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd123, 8'd45, 8'd32};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd120, 8'd41, 8'd26};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd122, 8'd43, 8'd28};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd128, 8'd47, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd115, 8'd34, 8'd17};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd115, 8'd38, 8'd20};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd117, 8'd41, 8'd27};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd113, 8'd41, 8'd27};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd88, 8'd18, 8'd8};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd94, 8'd24, 8'd14};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd126, 8'd54, 8'd40};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd126, 8'd50, 8'd36};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd118, 8'd41, 8'd23};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd124, 8'd43, 8'd26};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd115, 8'd34, 8'd17};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd109, 8'd30, 8'd13};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd115, 8'd36, 8'd19};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd117, 8'd40, 8'd22};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd110, 8'd35, 8'd16};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd107, 8'd32, 8'd13};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd108, 8'd33, 8'd14};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd98, 8'd27, 8'd5};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd96, 8'd31, 8'd9};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd89, 8'd32, 8'd12};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd61, 8'd9, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd66, 8'd14, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd97, 8'd40, 8'd20};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd100, 8'd35, 8'd13};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd94, 8'd23, 8'd1};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd85, 8'd20, 8'd16};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd79, 8'd22, 8'd13};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd77, 8'd25, 8'd12};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd83, 8'd27, 8'd14};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd92, 8'd25, 8'd17};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd88, 8'd20, 8'd17};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd70, 8'd15, 8'd12};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd52, 8'd11, 8'd5};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd68, 8'd20, 8'd6};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd105, 8'd47, 8'd33};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd111, 8'd39, 8'd24};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd105, 8'd29, 8'd15};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd94, 8'd26, 8'd17};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd69, 8'd19, 8'd20};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd99, 8'd72, 8'd81};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd123, 8'd112, 8'd128};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd100, 8'd119, 8'd134};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd61, 8'd88, 8'd83};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd61, 8'd91, 8'd93};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd74, 8'd93, 8'd126};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd104, 8'd104, 8'd130};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd180, 8'd160, 8'd127};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd240, 8'd195, 8'd110};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd91};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd131};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd101};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd244, 8'd215, 8'd77};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd240, 8'd224, 8'd89};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd245, 8'd237, 8'd136};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd249, 8'd251, 8'd188};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd252, 8'd227, 8'd186};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd235, 8'd195, 8'd126};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd224, 8'd174, 8'd75};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd221, 8'd153, 8'd42};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd64};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd255, 8'd142, 8'd59};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd223, 8'd74, 8'd42};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd242, 8'd58, 8'd50};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd248, 8'd51, 8'd61};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd229, 8'd59, 8'd62};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd222, 8'd61, 8'd53};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd234, 8'd55, 8'd50};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd240, 8'd52, 8'd53};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd58};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd215, 8'd39, 8'd39};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd213, 8'd37, 8'd37};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd213, 8'd34, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd184, 8'd35, 8'd3};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd229, 8'd111, 8'd39};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd244, 8'd138, 8'd29};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd239, 8'd130, 8'd13};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd236, 8'd134, 8'd34};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd189, 8'd114, 8'd49};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd221, 8'd172, 8'd132};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd115: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd205, 8'd147, 8'd109};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd221, 8'd111, 8'd32};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd115, 8'd10};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd237, 8'd143, 8'd21};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd47};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd214, 8'd92, 8'd19};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd177, 8'd33, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd192, 8'd28, 8'd26};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd212, 8'd34, 8'd46};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd219, 8'd33, 8'd46};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd231, 8'd44, 8'd53};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd237, 8'd52, 8'd57};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd242, 8'd58, 8'd68};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd237, 8'd57, 8'd68};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd224, 8'd57, 8'd48};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd233, 8'd92, 8'd47};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd62};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd253, 8'd169, 8'd53};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd217, 8'd148, 8'd18};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd240, 8'd214, 8'd153};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd246, 8'd229, 8'd186};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd251, 8'd236, 8'd171};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd240, 8'd214, 8'd127};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd253, 8'd196, 8'd80};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd90};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd94};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd81};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd64};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd243, 8'd161, 8'd59};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd217, 8'd163, 8'd73};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd198, 8'd169, 8'd89};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd116, 8'd132, 8'd122};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd83, 8'd93, 8'd94};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd95, 8'd102, 8'd112};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd99, 8'd109, 8'd121};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd102, 8'd117, 8'd124};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd82, 8'd91, 8'd86};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd66, 8'd54, 8'd40};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd57, 8'd26, 8'd6};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd75, 8'd28, 8'd20};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd84, 8'd28, 8'd13};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd88, 8'd25, 8'd7};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd86, 8'd27, 8'd13};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd94, 8'd45, 8'd40};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd56, 8'd11, 8'd8};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd100, 8'd47, 8'd41};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd103, 8'd41, 8'd28};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd95, 8'd35, 8'd25};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd77, 8'd17, 8'd6};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd103, 8'd43, 8'd32};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd100, 8'd38, 8'd25};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd97, 8'd34, 8'd19};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd98, 8'd35, 8'd20};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd105, 8'd39, 8'd23};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd93, 8'd27, 8'd11};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd99, 8'd36, 8'd19};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd98, 8'd36, 8'd21};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd95, 8'd37, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd73, 8'd19, 8'd7};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd78, 8'd24, 8'd12};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd106, 8'd48, 8'd36};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd105, 8'd43, 8'd28};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd99, 8'd36, 8'd19};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd106, 8'd38, 8'd25};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd96, 8'd28, 8'd15};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd91, 8'd25, 8'd11};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd97, 8'd31, 8'd17};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd98, 8'd35, 8'd20};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd92, 8'd30, 8'd15};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd88, 8'd26, 8'd11};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd87, 8'd28, 8'd12};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd81, 8'd20, 8'd17};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd77, 8'd21, 8'd20};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd71, 8'd23, 8'd23};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd48, 8'd4, 8'd5};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd52, 8'd8, 8'd9};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd79, 8'd31, 8'd31};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd80, 8'd24, 8'd23};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd77, 8'd16, 8'd13};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd68, 8'd17, 8'd13};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd62, 8'd19, 8'd10};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd59, 8'd21, 8'd8};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd67, 8'd23, 8'd10};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd75, 8'd22, 8'd14};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd72, 8'd17, 8'd14};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd53, 8'd12, 8'd8};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd37, 8'd8, 8'd4};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd46, 8'd10, 8'd0};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd87, 8'd41, 8'd26};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd97, 8'd41, 8'd26};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd92, 8'd30, 8'd17};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd81, 8'd26, 8'd19};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd61, 8'd22, 8'd27};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd109, 8'd91, 8'd105};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd109, 8'd104, 8'd126};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd111};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd47, 8'd58, 8'd62};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd64, 8'd70, 8'd84};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd77, 8'd67, 8'd104};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd121, 8'd89, 8'd104};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd200, 8'd147, 8'd95};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd235, 8'd158, 8'd54};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd45};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd255, 8'd186, 8'd70};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd78};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd78};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd66};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd66};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd252, 8'd214, 8'd105};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd176};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd253, 8'd234, 8'd191};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd238, 8'd201, 8'd123};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd218, 8'd155, 8'd58};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd249, 8'd160, 8'd60};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd255, 8'd153, 8'd60};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd228, 8'd87, 8'd44};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd239, 8'd59, 8'd45};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd245, 8'd49, 8'd59};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd233, 8'd60, 8'd64};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd223, 8'd60, 8'd55};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd235, 8'd53, 8'd49};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd241, 8'd53, 8'd54};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd228, 8'd53, 8'd58};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd44};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd214, 8'd38, 8'd38};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd211, 8'd35, 8'd35};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd218, 8'd36, 8'd33};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd179, 8'd20, 8'd1};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd199, 8'd65, 8'd14};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd252, 8'd133, 8'd43};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd246, 8'd132, 8'd17};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd238, 8'd133, 8'd24};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd203, 8'd118, 8'd38};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd201, 8'd131, 8'd82};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd116: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd225};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd182, 8'd111, 8'd57};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd243, 8'd126, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd118, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd241, 8'd144, 8'd27};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd252, 8'd141, 8'd51};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd177, 8'd46, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd184, 8'd31, 8'd13};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd198, 8'd28, 8'd29};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd207, 8'd27, 8'd36};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd217, 8'd33, 8'd43};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd231, 8'd46, 8'd54};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd239, 8'd53, 8'd58};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd247, 8'd62, 8'd76};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd235, 8'd59, 8'd70};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd224, 8'd67, 8'd50};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd243, 8'd113, 8'd51};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd63};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd247, 8'd167, 8'd54};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd217, 8'd150, 8'd35};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd242, 8'd237, 8'd207};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd241, 8'd218, 8'd142};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd243, 8'd199, 8'd76};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd249, 8'd190, 8'd36};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd49};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd253, 8'd189, 8'd40};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd247, 8'd176, 8'd26};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd249, 8'd164, 8'd11};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd252, 8'd158, 8'd10};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd246, 8'd159, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd227, 8'd163, 8'd63};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd213, 8'd167, 8'd90};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd100, 8'd122, 8'd119};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd60, 8'd73, 8'd79};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd69, 8'd75, 8'd91};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd65, 8'd73, 8'd92};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd76, 8'd92, 8'd107};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd62, 8'd75, 8'd81};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd59, 8'd58, 8'd54};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd54, 8'd39, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd61, 8'd31, 8'd7};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd67, 8'd30, 8'd1};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd74, 8'd30, 8'd0};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd66, 8'd25, 8'd0};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd77, 8'd45, 8'd24};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd48, 8'd19, 8'd3};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd86, 8'd50, 8'd28};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd85, 8'd41, 8'd14};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd78, 8'd38, 8'd13};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd58, 8'd18, 8'd0};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd84, 8'd42, 8'd17};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd78, 8'd37, 8'd9};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd74, 8'd30, 8'd1};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd77, 8'd32, 8'd3};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd83, 8'd38, 8'd7};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd71, 8'd26, 8'd0};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd85, 8'd40, 8'd7};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd81, 8'd37, 8'd8};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd79, 8'd40, 8'd11};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd60, 8'd24, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd65, 8'd29, 8'd3};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd87, 8'd48, 8'd19};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd84, 8'd40, 8'd11};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd81, 8'd36, 8'd3};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd89, 8'd39, 8'd12};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd79, 8'd29, 8'd2};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd73, 8'd26, 8'd0};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd79, 8'd32, 8'd4};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd81, 8'd36, 8'd7};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd75, 8'd31, 8'd2};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd71, 8'd27, 8'd0};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd71, 8'd30, 8'd0};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd66, 8'd21, 8'd0};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd58, 8'd20, 8'd1};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd55, 8'd22, 8'd5};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd35, 8'd8, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd40, 8'd13, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd63, 8'd30, 8'd13};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd61, 8'd23, 8'd4};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd62, 8'd17, 8'd0};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd54, 8'd19, 8'd0};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd47, 8'd21, 8'd0};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd45, 8'd24, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd51, 8'd26, 8'd0};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd60, 8'd24, 8'd0};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd56, 8'd20, 8'd0};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd39, 8'd14, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd22, 8'd10, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd0, 8'd0};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd58, 8'd28, 8'd0};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd69, 8'd33, 8'd1};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd67, 8'd26, 8'd0};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd62, 8'd26, 8'd2};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd50, 8'd28, 8'd14};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd99, 8'd94, 8'd91};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd89, 8'd94, 8'd98};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd64, 8'd81, 8'd89};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd47, 8'd64, 8'd58};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd83};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd80, 8'd72, 8'd85};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd129, 8'd105, 8'd81};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd207, 8'd167, 8'd72};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd225, 8'd166, 8'd28};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd244, 8'd171, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd211, 8'd168, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd229, 8'd175, 8'd14};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd248, 8'd183, 8'd31};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd252, 8'd183, 8'd27};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd245, 8'd181, 8'd23};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd242, 8'd186, 8'd47};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd250, 8'd202, 8'd102};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd151};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd237, 8'd239, 8'd218};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd252, 8'd218, 8'd157};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd216, 8'd158, 8'd74};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd238, 8'd158, 8'd61};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd66};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd231, 8'd100, 8'd48};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd235, 8'd60, 8'd41};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd242, 8'd48, 8'd56};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd236, 8'd63, 8'd69};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd224, 8'd59, 8'd57};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd235, 8'd51, 8'd49};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd241, 8'd53, 8'd54};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd227, 8'd53, 8'd55};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd44};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd214, 8'd38, 8'd38};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd211, 8'd35, 8'd35};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd212, 8'd33, 8'd29};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd184, 8'd17, 8'd11};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd171, 8'd23, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd245, 8'd117, 8'd46};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd251, 8'd137, 8'd23};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd232, 8'd128, 8'd7};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd220, 8'd125, 8'd33};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd192, 8'd103, 8'd43};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd242, 8'd218, 8'd208};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd117: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd233, 8'd193, 8'd158};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd187, 8'd103, 8'd33};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd245, 8'd129, 8'd18};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd255, 8'd127, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd247, 8'd140, 8'd34};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd231, 8'd110, 8'd37};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd161, 8'd18, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd197, 8'd35, 8'd33};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd202, 8'd27, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd206, 8'd27, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd212, 8'd34, 8'd34};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd52};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd236, 8'd50, 8'd51};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd246, 8'd62, 8'd74};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd229, 8'd58, 8'd66};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd224, 8'd74, 8'd49};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd250, 8'd128, 8'd53};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd58};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd236, 8'd162, 8'd55};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd223, 8'd157, 8'd61};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd241, 8'd227, 8'd182};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd231, 8'd199, 8'd114};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd242, 8'd192, 8'd69};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd55};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd227, 8'd198, 8'd58};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd220, 8'd194, 8'd57};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd215, 8'd187, 8'd52};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd218, 8'd179, 8'd48};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd226, 8'd175, 8'd58};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd233, 8'd179, 8'd91};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd231, 8'd188, 8'd137};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd227, 8'd195, 8'd172};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd143, 8'd154, 8'd156};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd77, 8'd77, 8'd89};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd56, 8'd47, 8'd68};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd48, 8'd39, 8'd66};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd71, 8'd72, 8'd93};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd69, 8'd71, 8'd86};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd60, 8'd53, 8'd61};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd46, 8'd27, 8'd33};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd54, 8'd24, 8'd24};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd62, 8'd23, 8'd16};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd68, 8'd21, 8'd11};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd60, 8'd17, 8'd11};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd67, 8'd32, 8'd36};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd50, 8'd19, 8'd25};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd76, 8'd40, 8'd42};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd76, 8'd31, 8'd26};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd71, 8'd33, 8'd32};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd51, 8'd11, 8'd11};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd74, 8'd34, 8'd32};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd67, 8'd26, 8'd24};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd61, 8'd20, 8'd16};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd65, 8'd22, 8'd16};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd72, 8'd29, 8'd23};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd62, 8'd17, 8'd11};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd77, 8'd33, 8'd24};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd70, 8'd27, 8'd20};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd69, 8'd30, 8'd25};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd54, 8'd19, 8'd17};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd58, 8'd23, 8'd21};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd75, 8'd36, 8'd31};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd71, 8'd28, 8'd21};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd69, 8'd25, 8'd16};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd79, 8'd30, 8'd26};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd69, 8'd20, 8'd16};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd64, 8'd16, 8'd12};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd70, 8'd22, 8'd18};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd71, 8'd26, 8'd21};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd65, 8'd22, 8'd16};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd61, 8'd18, 8'd12};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd62, 8'd19, 8'd13};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd62, 8'd17, 8'd0};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd52, 8'd14, 8'd0};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd49, 8'd18, 8'd0};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd33, 8'd7, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd38, 8'd12, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd57, 8'd26, 8'd8};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd55, 8'd17, 8'd0};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd58, 8'd13, 8'd0};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd50, 8'd14, 8'd16};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd44, 8'd16, 8'd13};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd39, 8'd19, 8'd10};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd47, 8'd20, 8'd13};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd56, 8'd18, 8'd15};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd53, 8'd14, 8'd15};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd34, 8'd8, 8'd11};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd16, 8'd4, 8'd4};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd20, 8'd0, 8'd0};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd48, 8'd17, 8'd15};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd58, 8'd19, 8'd12};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd59, 8'd19, 8'd9};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd57, 8'd22, 8'd16};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd57, 8'd32, 8'd35};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd86, 8'd75, 8'd89};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd77, 8'd75, 8'd96};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd40, 8'd61, 8'd88};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd24, 8'd46, 8'd60};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd43, 8'd59, 8'd75};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd68, 8'd73, 8'd95};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd149, 8'd146, 8'd131};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd233, 8'd224, 8'd149};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd239, 8'd216, 8'd122};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd246, 8'd213, 8'd134};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd222, 8'd216, 8'd94};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd224, 8'd214, 8'd80};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd228, 8'd209, 8'd70};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd233, 8'd203, 8'd83};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd237, 8'd200, 8'd111};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd242, 8'd205, 8'd134};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd244, 8'd217, 8'd140};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd247, 8'd226, 8'd135};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd205};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd175};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd217, 8'd158, 8'd82};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd232, 8'd158, 8'd61};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd69};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd236, 8'd112, 8'd52};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd230, 8'd60, 8'd35};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd240, 8'd47, 8'd52};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd239, 8'd64, 8'd71};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd226, 8'd58, 8'd58};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd234, 8'd50, 8'd50};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd242, 8'd54, 8'd55};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd225, 8'd53, 8'd53};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd216, 8'd40, 8'd40};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd214, 8'd38, 8'd38};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd210, 8'd34, 8'd34};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd202, 8'd27, 8'd22};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd187, 8'd16, 8'd22};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd158, 8'd1, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd224, 8'd89, 8'd34};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd252, 8'd138, 8'd26};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd229, 8'd128, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd226, 8'd128, 8'd19};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd202, 8'd98, 8'd27};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd215, 8'd186, 8'd172};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd118: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd198, 8'd139, 8'd97};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd205, 8'd109, 8'd33};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd238, 8'd124, 8'd12};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd248, 8'd134, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd249, 8'd135, 8'd39};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd198, 8'd67, 8'd11};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd171, 8'd18, 8'd10};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd201, 8'd31, 8'd44};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd201, 8'd24, 8'd32};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd211, 8'd37, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd208, 8'd37, 8'd27};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd218, 8'd49, 8'd44};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd235, 8'd48, 8'd43};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd240, 8'd59, 8'd68};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd223, 8'd54, 8'd59};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd223, 8'd78, 8'd47};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd251, 8'd136, 8'd53};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd248, 8'd161, 8'd48};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd229, 8'd155, 8'd56};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd234, 8'd167, 8'd89};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd161, 8'd156, 8'd118};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd97, 8'd78, 8'd48};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd73, 8'd40, 8'd21};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd68, 8'd36, 8'd23};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd87, 8'd64, 8'd48};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd87, 8'd71, 8'd46};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd71, 8'd50, 8'd21};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd56, 8'd25, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd58, 8'd19, 8'd4};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd68, 8'd20, 8'd0};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd69, 8'd13, 8'd0};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd66, 8'd14, 8'd0};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd66, 8'd22, 8'd11};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd62, 8'd22, 8'd14};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd79, 8'd33, 8'd20};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd80, 8'd25, 8'd5};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd79, 8'd33, 8'd17};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd58, 8'd11, 8'd0};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd80, 8'd33, 8'd17};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd72, 8'd23, 8'd6};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd65, 8'd17, 8'd0};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd70, 8'd19, 8'd0};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd78, 8'd26, 8'd5};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd68, 8'd16, 8'd0};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd80, 8'd26, 8'd2};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd70, 8'd20, 8'd0};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd69, 8'd22, 8'd2};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd59, 8'd14, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd62, 8'd17, 8'd0};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd74, 8'd27, 8'd7};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd68, 8'd18, 8'd0};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd71, 8'd17, 8'd0};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd80, 8'd21, 8'd3};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd69, 8'd12, 8'd0};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd65, 8'd8, 8'd0};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd70, 8'd15, 8'd0};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd71, 8'd19, 8'd0};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd66, 8'd14, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd61, 8'd10, 8'd0};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd62, 8'd11, 8'd0};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd71, 8'd12, 8'd6};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd60, 8'd7, 8'd1};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd58, 8'd10, 8'd6};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd45, 8'd4, 8'd2};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd50, 8'd9, 8'd7};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd67, 8'd19, 8'd15};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd63, 8'd10, 8'd4};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd67, 8'd8, 8'd2};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd60, 8'd14, 8'd0};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd53, 8'd16, 8'd0};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd51, 8'd19, 8'd0};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd57, 8'd21, 8'd0};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd66, 8'd19, 8'd1};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd62, 8'd14, 8'd0};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd45, 8'd9, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd27, 8'd5, 8'd0};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd50, 8'd13, 8'd4};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd67, 8'd25, 8'd9};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd67, 8'd21, 8'd0};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd74, 8'd24, 8'd0};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd72, 8'd28, 8'd1};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd77, 8'd45, 8'd24};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd79, 8'd57, 8'd44};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd79, 8'd66, 8'd60};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd76, 8'd71, 8'd77};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd63, 8'd58, 8'd54};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd71, 8'd65, 8'd65};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd107, 8'd97, 8'd106};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd190, 8'd181, 8'd166};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd252, 8'd245, 8'd193};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd254, 8'd241, 8'd199};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd193};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd219, 8'd159, 8'd87};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd229, 8'd154, 8'd52};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd252, 8'd176, 8'd56};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd239, 8'd120, 8'd54};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd226, 8'd61, 8'd31};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd236, 8'd46, 8'd48};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd240, 8'd64, 8'd74};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd227, 8'd58, 8'd61};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd235, 8'd49, 8'd50};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd243, 8'd55, 8'd56};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd223, 8'd54, 8'd51};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd216, 8'd40, 8'd40};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd213, 8'd37, 8'd37};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd211, 8'd35, 8'd35};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd210, 8'd34, 8'd34};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd195, 8'd24, 8'd17};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd185, 8'd13, 8'd25};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd164, 8'd0, 8'd9};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd194, 8'd55, 8'd14};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd246, 8'd136, 8'd25};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd232, 8'd137, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd221, 8'd121, 8'd1};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd221, 8'd108, 8'd28};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd187, 8'd154, 8'd137};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd119: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd181, 8'd110, 8'd66};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd216, 8'd112, 8'd39};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd231, 8'd120, 8'd15};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd242, 8'd139, 8'd10};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd251, 8'd129, 8'd43};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd172, 8'd35, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd189, 8'd31, 8'd32};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd197, 8'd24, 8'd44};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd199, 8'd22, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd217, 8'd45, 8'd33};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd205, 8'd38, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd211, 8'd49, 8'd38};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd222, 8'd45, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd223, 8'd44, 8'd47};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd56};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd54};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd232, 8'd55, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd234, 8'd56, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd234, 8'd54, 8'd63};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd239, 8'd52, 8'd43};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd244, 8'd63, 8'd68};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd225, 8'd59, 8'd63};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd230, 8'd88, 8'd52};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd255, 8'd148, 8'd59};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd250, 8'd164, 8'd51};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd232, 8'd159, 8'd64};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd248, 8'd180, 8'd115};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd232, 8'd215, 8'd127};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd211, 8'd198, 8'd93};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd213, 8'd195, 8'd97};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd186, 8'd152, 8'd63};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd194, 8'd147, 8'd69};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd198, 8'd150, 8'd78};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd192, 8'd154, 8'd79};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd185, 8'd156, 8'd76};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd183, 8'd151, 8'd66};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd193, 8'd153, 8'd66};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd188, 8'd148, 8'd52};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd199, 8'd150, 8'd47};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd197, 8'd140, 8'd33};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd197, 8'd144, 8'd42};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd192, 8'd149, 8'd55};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd196, 8'd156, 8'd68};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd206, 8'd160, 8'd66};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd208, 8'd153, 8'd53};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd213, 8'd167, 8'd71};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd191, 8'd145, 8'd49};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd212, 8'd166, 8'd68};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd204, 8'd156, 8'd56};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd198, 8'd148, 8'd49};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd201, 8'd152, 8'd50};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd210, 8'd158, 8'd57};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd200, 8'd148, 8'd46};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd207, 8'd154, 8'd48};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd198, 8'd147, 8'd42};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd197, 8'd149, 8'd47};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd187, 8'd141, 8'd43};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd190, 8'd144, 8'd46};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd202, 8'd154, 8'd52};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd195, 8'd144, 8'd39};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd196, 8'd143, 8'd37};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd207, 8'd149, 8'd50};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd197, 8'd139, 8'd40};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd191, 8'd136, 8'd36};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd197, 8'd142, 8'd42};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd199, 8'd145, 8'd45};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd193, 8'd141, 8'd40};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd189, 8'd137, 8'd36};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd190, 8'd138, 8'd37};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd205, 8'd149, 8'd38};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd193, 8'd142, 8'd33};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd191, 8'd147, 8'd40};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd181, 8'd143, 8'd36};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd186, 8'd148, 8'd41};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd200, 8'd156, 8'd49};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd196, 8'd145, 8'd36};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd201, 8'd145, 8'd34};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd194, 8'd148, 8'd52};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd188, 8'd150, 8'd49};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd185, 8'd154, 8'd48};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd192, 8'd155, 8'd49};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd201, 8'd153, 8'd53};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd197, 8'd148, 8'd53};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd179, 8'd143, 8'd47};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd162, 8'd139, 8'd43};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd172, 8'd135, 8'd46};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd183, 8'd140, 8'd45};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd177, 8'd130, 8'd26};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd183, 8'd135, 8'd24};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd182, 8'd139, 8'd26};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd191, 8'd159, 8'd50};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd171, 8'd149, 8'd48};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd179, 8'd164, 8'd69};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd197, 8'd158, 8'd81};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd195, 8'd157, 8'd72};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd194, 8'd156, 8'd83};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd197, 8'd161, 8'd103};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd218, 8'd188, 8'd118};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd221, 8'd197, 8'd111};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd219, 8'd194, 8'd138};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd212};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd225, 8'd162, 8'd93};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd228, 8'd147, 8'd40};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd248, 8'd167, 8'd36};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd242, 8'd125, 8'd55};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd225, 8'd62, 8'd29};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd235, 8'd45, 8'd47};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd241, 8'd65, 8'd75};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd228, 8'd58, 8'd61};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd235, 8'd49, 8'd50};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd244, 8'd56, 8'd57};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd223, 8'd54, 8'd51};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd216, 8'd40, 8'd40};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd213, 8'd37, 8'd37};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd211, 8'd35, 8'd35};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd210, 8'd34, 8'd34};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd191, 8'd24, 8'd16};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd181, 8'd9, 8'd25};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd173, 8'd8, 8'd25};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd172, 8'd32, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd240, 8'd132, 8'd21};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd237, 8'd146, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd215, 8'd113, 8'd0};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd239, 8'd121, 8'd34};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd169, 8'd134, 8'd115};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd120: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd251, 8'd198, 8'd164};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd195, 8'd86, 8'd17};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd244, 8'd129, 8'd23};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd232, 8'd127, 8'd12};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd243, 8'd136, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd212, 8'd69, 8'd37};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd180, 8'd28, 8'd5};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd174, 8'd7, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd204, 8'd25, 8'd28};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd218, 8'd37, 8'd44};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd205, 8'd28, 8'd34};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd204, 8'd36, 8'd35};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd219, 8'd57, 8'd52};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd44};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd229, 8'd53, 8'd53};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd231, 8'd55, 8'd55};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd231, 8'd55, 8'd55};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd228, 8'd65, 8'd56};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd232, 8'd49, 8'd54};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd221, 8'd58, 8'd51};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd201, 8'd88, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd59};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd248, 8'd150, 8'd43};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd214, 8'd143, 8'd65};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd235, 8'd214, 8'd161};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd232, 8'd194, 8'd113};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd220, 8'd148, 8'd38};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd255, 8'd170, 8'd52};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd249, 8'd197, 8'd75};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd253, 8'd198, 8'd81};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd83};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd252, 8'd189, 8'd84};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd252, 8'd187, 8'd85};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd254, 8'd191, 8'd88};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd91};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd92};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd85};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd250, 8'd196, 8'd70};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd71};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd249, 8'd192, 8'd61};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd74};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd243, 8'd195, 8'd69};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd86};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd245, 8'd210, 8'd94};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd80};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd250, 8'd214, 8'd91};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd102};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd102};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd90};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd253, 8'd194, 8'd76};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd66};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd61};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd250, 8'd196, 8'd70};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd239, 8'd185, 8'd61};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd245, 8'd189, 8'd68};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd86};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd83};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd238, 8'd176, 8'd65};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd237, 8'd175, 8'd66};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd84};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd246, 8'd181, 8'd65};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd242, 8'd179, 8'd63};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd239, 8'd176, 8'd60};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd235, 8'd174, 8'd57};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd233, 8'd174, 8'd56};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd233, 8'd177, 8'd58};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd234, 8'd179, 8'd60};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd233, 8'd181, 8'd61};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd243, 8'd187, 8'd38};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd244, 8'd187, 8'd46};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd247, 8'd187, 8'd57};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd246, 8'd186, 8'd64};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd244, 8'd185, 8'd65};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd239, 8'd186, 8'd58};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd233, 8'd186, 8'd46};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd230, 8'd186, 8'd38};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd226, 8'd176, 8'd65};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd72};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd239, 8'd191, 8'd80};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd238, 8'd192, 8'd80};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd225, 8'd182, 8'd69};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd217, 8'd174, 8'd61};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd224, 8'd183, 8'd69};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd239, 8'd198, 8'd84};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd247, 8'd183, 8'd73};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd233, 8'd171, 8'd60};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd222, 8'd166, 8'd57};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd224, 8'd173, 8'd68};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd227, 8'd182, 8'd79};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd224, 8'd185, 8'd84};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd222, 8'd186, 8'd89};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd224, 8'd190, 8'd93};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd223, 8'd186, 8'd105};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd241, 8'd214, 8'd133};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd233, 8'd212, 8'd133};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd245, 8'd216, 8'd140};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd247, 8'd201, 8'd124};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd225, 8'd167, 8'd85};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd203, 8'd147, 8'd52};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd241, 8'd189, 8'd87};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd246, 8'd213, 8'd172};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd218, 8'd147, 8'd57};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd253, 8'd155, 8'd28};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd255, 8'd162, 8'd56};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd216, 8'd83, 8'd52};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd219, 8'd58, 8'd73};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd229, 8'd56, 8'd52};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd237, 8'd55, 8'd41};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd231, 8'd48, 8'd50};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd238, 8'd64, 8'd65};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd213, 8'd49, 8'd22};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd228, 8'd50, 8'd50};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd228, 8'd50, 8'd50};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd216, 8'd42, 8'd41};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd210, 8'd36, 8'd35};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd203, 8'd31, 8'd29};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd200, 8'd28, 8'd26};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd181, 8'd19, 8'd0};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd184, 8'd10, 8'd12};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd177, 8'd0, 8'd13};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd160, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd223, 8'd93, 8'd31};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd243, 8'd138, 8'd31};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd222, 8'd124, 8'd1};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd225, 8'd125, 8'd3};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd177, 8'd87, 8'd9};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd171};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd121: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd219, 8'd163, 8'd126};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd215, 8'd105, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd239, 8'd124, 8'd17};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd233, 8'd128, 8'd13};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd246, 8'd137, 8'd34};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd196, 8'd51, 8'd22};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd174, 8'd19, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd171, 8'd4, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd195, 8'd19, 8'd21};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd211, 8'd30, 8'd35};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd204, 8'd28, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd201, 8'd33, 8'd32};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd212, 8'd49, 8'd44};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd44};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd229, 8'd53, 8'd53};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd231, 8'd55, 8'd55};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd234, 8'd65, 8'd58};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd236, 8'd51, 8'd56};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd219, 8'd57, 8'd46};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd225, 8'd111, 8'd49};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd254, 8'd161, 8'd58};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd246, 8'd153, 8'd50};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd221, 8'd154, 8'd83};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd245, 8'd227, 8'd179};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd232};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd236, 8'd211, 8'd144};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd218, 8'd170, 8'd62};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd235, 8'd157, 8'd31};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd253, 8'd158, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd249, 8'd178, 8'd64};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd245, 8'd171, 8'd62};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd248, 8'd171, 8'd67};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd79};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd255, 8'd174, 8'd80};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd249, 8'd166, 8'd70};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd249, 8'd167, 8'd68};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd75};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd251, 8'd172, 8'd69};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd251, 8'd168, 8'd64};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd253, 8'd166, 8'd60};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd251, 8'd163, 8'd55};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd72};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd81};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd89};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd248, 8'd175, 8'd81};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd251, 8'd194, 8'd87};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd254, 8'd192, 8'd89};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd255, 8'd188, 8'd89};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd255, 8'd181, 8'd84};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd176, 8'd77};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd255, 8'd177, 8'd72};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd69};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd68};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd69};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd255, 8'd184, 8'd68};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd72};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd76};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd255, 8'd180, 8'd74};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd250, 8'd171, 8'd68};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd72};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd82};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd249, 8'd186, 8'd81};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd250, 8'd187, 8'd82};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd250, 8'd189, 8'd83};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd248, 8'd191, 8'd84};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd247, 8'd193, 8'd85};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd246, 8'd195, 8'd86};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd244, 8'd196, 8'd86};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd244, 8'd196, 8'd86};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd80};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd84};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd89};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd92};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd91};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd88};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd83};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd78};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd104};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd106};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd108};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd107};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd101};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd255, 8'd192, 8'd98};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd100};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd104};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd102};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd255, 8'd187, 8'd90};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd248, 8'd182, 8'd88};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd103};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd119};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd126};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd125};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd211, 8'd126};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd141};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd160};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd161};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd169};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd153};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd250, 8'd191, 8'd113};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd218, 8'd162, 8'd69};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd227, 8'd178, 8'd75};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd244, 8'd212, 8'd173};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd218};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd251, 8'd221, 8'd183};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd227, 8'd161, 8'd77};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd244, 8'd151, 8'd32};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd255, 8'd156, 8'd47};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd232, 8'd105, 8'd62};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd214, 8'd60, 8'd60};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd228, 8'd57, 8'd49};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd232, 8'd52, 8'd38};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd236, 8'd53, 8'd57};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd235, 8'd59, 8'd62};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd218, 8'd51, 8'd32};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd227, 8'd49, 8'd49};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd227, 8'd49, 8'd49};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd215, 8'd41, 8'd40};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd209, 8'd35, 8'd34};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd202, 8'd30, 8'd28};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd198, 8'd26, 8'd24};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd180, 8'd19, 8'd0};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd183, 8'd11, 8'd11};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd176, 8'd0, 8'd12};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd160, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd207, 8'd77, 8'd19};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd241, 8'd133, 8'd32};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd228, 8'd129, 8'd9};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd228, 8'd125, 8'd4};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd188, 8'd97, 8'd18};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd242, 8'd190, 8'd142};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd122: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd184, 8'd121, 8'd77};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd233, 8'd123, 8'd38};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd231, 8'd121, 8'd6};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd237, 8'd132, 8'd17};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd244, 8'd131, 8'd35};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd176, 8'd27, 8'd3};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd166, 8'd11, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd168, 8'd1, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd185, 8'd11, 8'd10};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd202, 8'd23, 8'd27};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd203, 8'd27, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd201, 8'd31, 8'd31};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd203, 8'd38, 8'd36};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd228, 8'd52, 8'd52};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd231, 8'd55, 8'd55};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd240, 8'd60, 8'd59};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd237, 8'd53, 8'd53};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd220, 8'd61, 8'd39};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd138, 8'd71};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd252, 8'd158, 8'd58};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd237, 8'd153, 8'd57};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd230, 8'd176, 8'd112};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd206};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd255, 8'd221};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd247, 8'd221, 8'd146};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd216, 8'd171, 8'd54};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd221, 8'd154, 8'd13};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd241, 8'd154, 8'd13};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd243, 8'd142, 8'd10};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd210, 8'd108, 8'd8};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd193, 8'd91, 8'd0};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd189, 8'd86, 8'd0};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd202, 8'd96, 8'd10};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd201, 8'd95, 8'd9};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd191, 8'd82, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd194, 8'd84, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd209, 8'd100, 8'd9};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd199, 8'd82, 8'd3};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd202, 8'd83, 8'd3};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd202, 8'd79, 8'd0};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd214, 8'd89, 8'd7};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd219, 8'd94, 8'd14};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd227, 8'd105, 8'd28};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd221, 8'd100, 8'd27};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd216, 8'd99, 8'd29};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd199, 8'd106, 8'd26};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd200, 8'd104, 8'd20};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd202, 8'd102, 8'd14};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd206, 8'd101, 8'd9};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd212, 8'd103, 8'd10};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd211, 8'd104, 8'd10};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd209, 8'd101, 8'd10};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd204, 8'd99, 8'd8};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd194, 8'd97, 8'd0};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd203, 8'd106, 8'd3};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd208, 8'd109, 8'd8};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd204, 8'd104, 8'd6};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd200, 8'd97, 8'd4};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd199, 8'd94, 8'd3};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd197, 8'd91, 8'd3};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd195, 8'd89, 8'd1};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd213, 8'd96, 8'd19};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd210, 8'd94, 8'd17};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd204, 8'd91, 8'd13};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd199, 8'd89, 8'd10};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd195, 8'd90, 8'd9};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd192, 8'd91, 8'd9};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd194, 8'd95, 8'd12};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd193, 8'd97, 8'd13};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd191, 8'd102, 8'd8};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd195, 8'd105, 8'd17};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd199, 8'd110, 8'd28};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd202, 8'd112, 8'd36};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd200, 8'd113, 8'd36};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd195, 8'd110, 8'd27};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd190, 8'd106, 8'd16};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd186, 8'd103, 8'd7};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd197, 8'd107, 8'd29};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd198, 8'd108, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd198, 8'd106, 8'd29};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd198, 8'd106, 8'd29};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd203, 8'd110, 8'd33};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd208, 8'd115, 8'd38};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd209, 8'd113, 8'd37};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd204, 8'd108, 8'd32};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd189, 8'd100, 8'd20};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd184, 8'd97, 8'd17};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd187, 8'd102, 8'd22};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd196, 8'd114, 8'd38};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd200, 8'd122, 8'd47};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd196, 8'd122, 8'd47};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd194, 8'd125, 8'd50};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd198, 8'd130, 8'd57};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd222, 8'd151, 8'd99};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd219, 8'd160, 8'd104};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd212, 8'd163, 8'd105};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd231, 8'd179, 8'd119};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd235, 8'd172, 8'd105};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd234, 8'd165, 8'd87};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd208, 8'd145, 8'd50};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd196, 8'd142, 8'd36};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd217, 8'd164, 8'd86};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd247, 8'd215, 8'd168};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd239, 8'd183, 8'd109};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd229, 8'd148, 8'd43};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd248, 8'd148, 8'd37};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd135, 8'd74};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd213, 8'd68, 8'd47};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd221, 8'd58, 8'd43};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd226, 8'd49, 8'd39};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd236, 8'd55, 8'd60};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd231, 8'd54, 8'd60};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd226, 8'd55, 8'd47};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd227, 8'd49, 8'd49};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd226, 8'd48, 8'd48};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd213, 8'd39, 8'd38};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd206, 8'd32, 8'd31};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd198, 8'd26, 8'd24};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd195, 8'd23, 8'd21};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd180, 8'd21, 8'd2};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd184, 8'd12, 8'd12};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd173, 8'd0, 8'd8};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd161, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd182, 8'd47, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd234, 8'd125, 8'd34};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd239, 8'd138, 8'd22};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd229, 8'd125, 8'd2};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd208, 8'd112, 8'd28};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd207, 8'd150, 8'd97};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd123: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd242, 8'd230, 8'd208};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd172, 8'd99, 8'd44};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd234, 8'd124, 8'd27};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd230, 8'd124, 8'd2};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd244, 8'd140, 8'd29};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd231, 8'd112, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd161, 8'd9, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd162, 8'd4, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd167, 8'd2, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd180, 8'd8, 8'd6};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd193, 8'd19, 8'd20};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd204, 8'd30, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd204, 8'd34, 8'd34};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd201, 8'd33, 8'd32};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd228, 8'd52, 8'd52};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd54};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd54};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd243, 8'd54, 8'd58};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd229, 8'd52, 8'd44};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd225, 8'd76, 8'd36};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd75};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd251, 8'd157, 8'd61};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd222, 8'd150, 8'd65};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd241, 8'd202, 8'd147};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd167};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd215, 8'd168, 8'd50};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd224, 8'd154, 8'd6};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd1};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd238, 8'd136, 8'd0};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd232, 8'd124, 8'd0};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd234, 8'd106, 8'd19};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd219, 8'd90, 8'd7};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd212, 8'd85, 8'd6};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd220, 8'd93, 8'd16};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd222, 8'd95, 8'd18};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd216, 8'd85, 8'd7};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd219, 8'd83, 8'd5};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd228, 8'd91, 8'd10};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd227, 8'd90, 8'd18};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd227, 8'd89, 8'd17};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd224, 8'd83, 8'd12};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd243, 8'd102, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd236, 8'd93, 8'd23};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd244, 8'd101, 8'd31};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd242, 8'd101, 8'd32};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd255, 8'd115, 8'd49};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd226, 8'd103, 8'd35};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd221, 8'd98, 8'd21};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd222, 8'd94, 8'd5};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd225, 8'd97, 8'd0};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd232, 8'd102, 8'd4};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd234, 8'd105, 8'd13};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd229, 8'd100, 8'd17};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd220, 8'd94, 8'd17};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd220, 8'd101, 8'd9};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd227, 8'd108, 8'd16};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd231, 8'd112, 8'd22};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd226, 8'd104, 8'd19};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd222, 8'd97, 8'd15};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd219, 8'd94, 8'd14};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd219, 8'd92, 8'd15};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd217, 8'd89, 8'd14};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd232, 8'd78, 8'd14};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd231, 8'd79, 8'd14};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd228, 8'd79, 8'd13};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd225, 8'd80, 8'd13};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd226, 8'd85, 8'd16};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd227, 8'd90, 8'd20};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd228, 8'd94, 8'd23};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd230, 8'd98, 8'd26};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd222, 8'd106, 8'd21};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd219, 8'd104, 8'd21};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd216, 8'd103, 8'd25};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd214, 8'd102, 8'd26};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd213, 8'd103, 8'd24};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd216, 8'd105, 8'd23};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd219, 8'd108, 8'd19};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd223, 8'd110, 8'd18};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd218, 8'd107, 8'd36};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd219, 8'd108, 8'd37};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd218, 8'd105, 8'd35};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd214, 8'd100, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd217, 8'd100, 8'd31};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd222, 8'd103, 8'd35};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd219, 8'd100, 8'd32};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd214, 8'd92, 8'd25};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd198, 8'd86, 8'd14};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd195, 8'd84, 8'd12};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd201, 8'd90, 8'd19};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd211, 8'd104, 8'd32};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd214, 8'd110, 8'd39};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd210, 8'd108, 8'd36};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd207, 8'd106, 8'd34};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd211, 8'd110, 8'd40};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd212, 8'd107, 8'd59};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd203, 8'd113, 8'd61};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd201, 8'd124, 8'd68};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd223, 8'd145, 8'd83};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd223, 8'd139, 8'd69};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd243, 8'd154, 8'd70};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd233, 8'd151, 8'd49};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd212, 8'd141, 8'd25};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd209, 8'd133, 8'd21};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd230, 8'd171, 8'd103};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd211};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd251, 8'd206, 8'd147};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd218, 8'd150, 8'd65};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd237, 8'd143, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd77};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd222, 8'd90, 8'd42};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd212, 8'd58, 8'd34};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd227, 8'd56, 8'd48};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd232, 8'd53, 8'd59};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd232, 8'd53, 8'd59};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd231, 8'd55, 8'd57};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd226, 8'd48, 8'd48};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd225, 8'd47, 8'd47};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd221, 8'd45, 8'd45};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd210, 8'd36, 8'd35};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd202, 8'd28, 8'd27};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd194, 8'd22, 8'd20};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd190, 8'd18, 8'd16};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd176, 8'd18, 8'd6};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd181, 8'd11, 8'd11};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd172, 8'd0, 8'd4};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd162, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd157, 8'd20, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd224, 8'd111, 8'd35};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd249, 8'd144, 8'd35};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd232, 8'd127, 8'd2};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd228, 8'd127, 8'd35};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd176, 8'd114, 8'd55};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd124: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd227, 8'd202, 8'd172};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd186, 8'd103, 8'd35};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd226, 8'd116, 8'd5};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd234, 8'd132, 8'd4};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd250, 8'd144, 8'd44};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd208, 8'd80, 8'd17};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd158, 8'd1, 8'd0};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd163, 8'd4, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd169, 8'd6, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd176, 8'd7, 8'd2};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd190, 8'd18, 8'd16};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd203, 8'd31, 8'd31};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd208, 8'd35, 8'd37};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd205, 8'd32, 8'd34};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd44};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd223, 8'd47, 8'd47};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd227, 8'd51, 8'd51};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd229, 8'd53, 8'd53};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd54};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd237, 8'd48, 8'd54};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd219, 8'd57, 8'd36};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd234, 8'd101, 8'd44};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd63};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd247, 8'd157, 8'd61};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd211, 8'd154, 8'd77};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd248, 8'd223, 8'd182};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd214};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd237, 8'd196, 8'd106};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd214, 8'd146, 8'd9};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd239, 8'd148, 8'd0};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd9};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd241, 8'd127, 8'd5};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd223, 8'd106, 8'd1};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd241, 8'd98, 8'd22};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd234, 8'd94, 8'd19};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd228, 8'd91, 8'd19};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd229, 8'd95, 8'd24};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd236, 8'd99, 8'd29};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd239, 8'd98, 8'd26};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd238, 8'd92, 8'd17};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd236, 8'd86, 8'd10};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd233, 8'd95, 8'd20};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd230, 8'd92, 8'd17};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd216, 8'd80, 8'd4};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd225, 8'd92, 8'd17};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd221, 8'd88, 8'd11};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd237, 8'd104, 8'd27};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd237, 8'd101, 8'd23};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd245, 8'd110, 8'd29};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd252, 8'd116, 8'd42};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd245, 8'd108, 8'd27};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd239, 8'd102, 8'd8};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd239, 8'd102, 8'd0};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd244, 8'd107, 8'd3};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd245, 8'd111, 8'd14};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd241, 8'd110, 8'd22};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd235, 8'd106, 8'd25};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd236, 8'd110, 8'd26};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd235, 8'd109, 8'd25};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd237, 8'd108, 8'd27};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd235, 8'd104, 8'd26};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd228, 8'd96, 8'd22};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd222, 8'd88, 8'd17};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd224, 8'd89, 8'd21};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd232, 8'd94, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd220, 8'd93, 8'd12};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd221, 8'd94, 8'd13};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd222, 8'd97, 8'd15};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd221, 8'd99, 8'd16};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd221, 8'd100, 8'd17};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd221, 8'd100, 8'd17};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd219, 8'd100, 8'd16};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd219, 8'd100, 8'd16};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd234, 8'd99, 8'd7};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd232, 8'd101, 8'd10};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd232, 8'd105, 8'd12};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd231, 8'd108, 8'd14};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd233, 8'd109, 8'd13};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd235, 8'd108, 8'd11};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd239, 8'd107, 8'd7};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd242, 8'd106, 8'd4};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd222, 8'd102, 8'd26};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd225, 8'd105, 8'd29};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd228, 8'd106, 8'd31};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd227, 8'd105, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd227, 8'd103, 8'd29};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd228, 8'd104, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd230, 8'd106, 8'd32};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd234, 8'd108, 8'd34};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd220, 8'd94, 8'd20};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd213, 8'd87, 8'd13};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd215, 8'd89, 8'd15};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd227, 8'd101, 8'd25};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd235, 8'd109, 8'd33};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd230, 8'd104, 8'd27};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd225, 8'd99, 8'd22};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd223, 8'd97, 8'd20};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd222, 8'd93, 8'd38};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd212, 8'd96, 8'd39};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd211, 8'd109, 8'd45};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd224, 8'd123, 8'd55};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd211, 8'd104, 8'd26};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd231, 8'd120, 8'd28};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd232, 8'd130, 8'd20};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd219, 8'd127, 8'd4};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd216, 8'd128, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd211, 8'd135, 8'd41};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd238, 8'd184, 8'd138};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd184};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd217, 8'd164, 8'd98};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd231, 8'd143, 8'd35};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd166, 8'd65};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd240, 8'd119, 8'd46};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd208, 8'd64, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd228, 8'd63, 8'd59};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd224, 8'd50, 8'd52};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd233, 8'd54, 8'd58};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd234, 8'd53, 8'd60};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd225, 8'd47, 8'd47};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd224, 8'd46, 8'd46};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd214, 8'd38, 8'd38};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd206, 8'd32, 8'd31};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd198, 8'd24, 8'd23};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd190, 8'd18, 8'd16};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd185, 8'd13, 8'd11};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd173, 8'd16, 8'd7};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd177, 8'd9, 8'd8};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd171, 8'd0, 8'd2};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd161, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd142, 8'd4, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd209, 8'd94, 8'd31};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd253, 8'd145, 8'd44};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd237, 8'd129, 8'd3};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd243, 8'd135, 8'd37};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd165, 8'd97, 8'd32};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd253, 8'd233, 8'd209};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd125: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd210, 8'd175, 8'd137};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd207, 8'd116, 8'd35};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd224, 8'd114, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd239, 8'd140, 8'd11};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd244, 8'd136, 8'd46};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd183, 8'd47, 8'd5};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd161, 8'd1, 8'd1};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd166, 8'd4, 8'd2};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd169, 8'd6, 8'd1};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd172, 8'd7, 8'd1};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd184, 8'd15, 8'd10};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd199, 8'd27, 8'd25};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd208, 8'd34, 8'd36};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd210, 8'd35, 8'd40};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd220, 8'd44, 8'd44};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd225, 8'd49, 8'd49};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd227, 8'd51, 8'd51};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd229, 8'd53, 8'd53};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd230, 8'd54, 8'd54};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd230, 8'd47, 8'd52};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd215, 8'd72, 8'd38};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd243, 8'd130, 8'd52};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd49};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd241, 8'd154, 8'd61};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd216, 8'd173, 8'd105};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd226, 8'd184, 8'd124};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd221, 8'd161, 8'd49};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd240, 8'd159, 8'd16};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd241, 8'd138, 8'd0};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd248, 8'd132, 8'd11};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd248, 8'd126, 8'd25};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd219, 8'd96, 8'd3};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd236, 8'd94, 8'd22};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd224, 8'd87, 8'd15};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd209, 8'd78, 8'd8};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd202, 8'd75, 8'd4};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd212, 8'd84, 8'd13};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd228, 8'd94, 8'd21};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd235, 8'd93, 8'd17};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd234, 8'd87, 8'd10};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd235, 8'd102, 8'd25};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd230, 8'd100, 8'd24};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd213, 8'd90, 8'd13};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd211, 8'd91, 8'd15};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd217, 8'd102, 8'd22};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd237, 8'd122, 8'd39};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd234, 8'd118, 8'd31};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd223, 8'd108, 8'd17};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd237, 8'd107, 8'd21};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd237, 8'd107, 8'd19};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd239, 8'd109, 8'd15};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd240, 8'd110, 8'd14};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd239, 8'd111, 8'd14};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd231, 8'd108, 8'd12};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd220, 8'd103, 8'd10};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd211, 8'd98, 8'd6};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd219, 8'd98, 8'd17};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd223, 8'd102, 8'd23};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd229, 8'd107, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd233, 8'd109, 8'd35};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd227, 8'd100, 8'd29};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd214, 8'd87, 8'd20};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd208, 8'd79, 8'd14};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd209, 8'd80, 8'd15};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd222, 8'd101, 8'd18};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd218, 8'd97, 8'd14};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd214, 8'd92, 8'd9};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd211, 8'd89, 8'd6};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd215, 8'd90, 8'd8};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd222, 8'd95, 8'd14};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd232, 8'd103, 8'd22};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd237, 8'd108, 8'd27};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd227, 8'd94, 8'd1};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd226, 8'd98, 8'd1};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd225, 8'd103, 8'd4};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd225, 8'd108, 8'd5};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd228, 8'd110, 8'd4};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd234, 8'd109, 8'd3};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd238, 8'd105, 8'd0};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd242, 8'd103, 8'd0};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd230, 8'd110, 8'd32};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd225, 8'd105, 8'd27};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd227, 8'd107, 8'd29};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd232, 8'd115, 8'd36};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd228, 8'd113, 8'd33};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd218, 8'd105, 8'd25};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd220, 8'd107, 8'd27};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd229, 8'd118, 8'd37};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd219, 8'd97, 8'd24};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd223, 8'd101, 8'd26};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd232, 8'd109, 8'd32};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd237, 8'd114, 8'd36};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd232, 8'd107, 8'd25};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd224, 8'd98, 8'd14};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd229, 8'd103, 8'd18};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd244, 8'd115, 8'd31};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd239, 8'd103, 8'd41};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd222, 8'd100, 8'd35};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd209, 8'd100, 8'd33};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd213, 8'd105, 8'd33};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd197, 8'd80, 8'd1};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd217, 8'd96, 8'd5};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd233, 8'd121, 8'd13};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd242, 8'd138, 8'd17};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd224, 8'd134, 8'd0};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd209, 8'd122, 8'd6};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd221, 8'd147, 8'd60};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd248, 8'd201, 8'd147};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd251, 8'd237, 8'd208};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd224, 8'd186, 8'd139};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd230, 8'd146, 8'd47};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd252, 8'd161, 8'd47};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd255, 8'd146, 8'd51};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd218, 8'd81, 8'd39};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd224, 8'd65, 8'd61};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd222, 8'd50, 8'd48};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd232, 8'd53, 8'd49};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd235, 8'd50, 8'd56};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd224, 8'd46, 8'd46};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd222, 8'd44, 8'd44};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd212, 8'd36, 8'd36};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd203, 8'd29, 8'd28};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd195, 8'd21, 8'd20};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd186, 8'd14, 8'd12};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd181, 8'd9, 8'd7};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd166, 8'd11, 8'd6};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd170, 8'd5, 8'd1};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd169, 8'd0, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd160, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd138, 8'd0, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd193, 8'd72, 8'd25};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd253, 8'd143, 8'd48};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd242, 8'd133, 8'd6};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd250, 8'd134, 8'd31};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd175, 8'd101, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd235, 8'd210, 8'd180};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd126: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd200, 8'd156, 8'd109};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd220, 8'd122, 8'd31};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd237, 8'd125, 8'd0};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd242, 8'd145, 8'd15};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd230, 8'd120, 8'd43};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd163, 8'd21, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd167, 8'd4, 8'd9};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd165, 8'd2, 8'd5};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd164, 8'd2, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd168, 8'd5, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd177, 8'd10, 8'd2};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd187, 8'd18, 8'd15};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd203, 8'd29, 8'd31};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd213, 8'd36, 8'd44};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd218, 8'd42, 8'd42};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd227, 8'd51, 8'd51};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd228, 8'd52, 8'd52};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd229, 8'd53, 8'd53};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd222, 8'd49, 8'd51};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd220, 8'd97, 8'd53};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd250, 8'd155, 8'd61};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd249, 8'd148, 8'd42};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd230, 8'd147, 8'd55};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd234, 8'd202, 8'd141};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd137};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd214, 8'd150, 8'd52};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd223, 8'd149, 8'd14};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd250, 8'd162, 8'd13};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd236, 8'd132, 8'd1};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd234, 8'd116, 8'd10};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd241, 8'd116, 8'd24};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd226, 8'd98, 8'd7};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd225, 8'd93, 8'd21};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd80, 8'd9};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd193, 8'd75, 8'd3};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd197, 8'd85, 8'd11};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd210, 8'd97, 8'd21};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd222, 8'd100, 8'd23};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd228, 8'd97, 8'd17};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd231, 8'd94, 8'd14};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd202, 8'd67, 8'd3};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd194, 8'd65, 8'd0};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd198, 8'd78, 8'd15};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd202, 8'd93, 8'd28};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd205, 8'd103, 8'd31};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd193, 8'd93, 8'd17};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd198, 8'd98, 8'd13};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd206, 8'd106, 8'd18};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd226, 8'd111, 8'd20};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd228, 8'd112, 8'd25};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd230, 8'd111, 8'd31};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd224, 8'd107, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd214, 8'd101, 8'd23};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd204, 8'd97, 8'd15};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd196, 8'd98, 8'd9};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd193, 8'd100, 8'd5};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd190, 8'd83, 8'd1};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd201, 8'd94, 8'd14};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd204, 8'd97, 8'd19};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd197, 8'd87, 8'd12};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd190, 8'd78, 8'd6};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd187, 8'd74, 8'd6};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd184, 8'd69, 8'd4};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd178, 8'd63, 8'd0};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd191, 8'd78, 8'd2};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd193, 8'd77, 8'd2};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd197, 8'd76, 8'd3};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd202, 8'd78, 8'd6};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd213, 8'd82, 8'd12};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd226, 8'd89, 8'd21};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd235, 8'd96, 8'd29};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd242, 8'd100, 8'd34};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd209, 8'd94, 8'd14};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd201, 8'd92, 8'd9};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd191, 8'd90, 8'd0};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd184, 8'd90, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd189, 8'd93, 8'd0};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd203, 8'd96, 8'd0};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd218, 8'd101, 8'd6};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd228, 8'd105, 8'd11};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd233, 8'd116, 8'd47};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd209, 8'd95, 8'd25};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd202, 8'd91, 8'd20};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd214, 8'd107, 8'd35};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd211, 8'd109, 8'd35};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd190, 8'd92, 8'd17};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd182, 8'd89, 8'd12};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd192, 8'd100, 8'd23};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd189, 8'd91, 8'd20};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd192, 8'd91, 8'd19};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd198, 8'd96, 8'd22};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd203, 8'd100, 8'd23};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd203, 8'd96, 8'd16};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd201, 8'd92, 8'd9};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd210, 8'd100, 8'd13};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd225, 8'd113, 8'd27};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd217, 8'd95, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd201, 8'd92, 8'd27};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd190, 8'd93, 8'd25};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd203, 8'd104, 8'd36};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd195, 8'd84, 8'd13};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd206, 8'd91, 8'd10};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd217, 8'd107, 8'd12};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd235, 8'd134, 8'd28};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd219, 8'd134, 8'd5};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd225, 8'd133, 8'd0};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd221, 8'd132, 8'd4};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd220, 8'd155, 8'd65};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd238, 8'd206, 8'd168};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd237, 8'd208, 8'd176};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd231, 8'd150, 8'd59};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd236, 8'd152, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd56};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd238, 8'd107, 8'd61};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd213, 8'd58, 8'd54};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd225, 8'd56, 8'd49};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd228, 8'd50, 8'd38};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd234, 8'd48, 8'd53};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd223, 8'd45, 8'd45};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd221, 8'd43, 8'd43};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd216, 8'd40, 8'd40};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd210, 8'd34, 8'd34};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd201, 8'd27, 8'd26};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd192, 8'd18, 8'd17};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd183, 8'd11, 8'd9};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd178, 8'd6, 8'd4};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd161, 8'd7, 8'd5};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd165, 8'd2, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd170, 8'd1, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd159, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd143, 8'd1, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd179, 8'd55, 8'd19};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd250, 8'd136, 8'd48};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd248, 8'd136, 8'd8};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd249, 8'd131, 8'd21};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd194, 8'd116, 8'd41};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd215, 8'd189, 8'd156};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd127: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd197, 8'd147, 8'd94};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd221, 8'd121, 8'd25};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd252, 8'd139, 8'd7};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd240, 8'd145, 8'd17};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd214, 8'd106, 8'd34};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd155, 8'd8, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd170, 8'd4, 8'd14};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd163, 8'd0, 8'd3};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd160, 8'd0, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd165, 8'd2, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd170, 8'd6, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd180, 8'd11, 8'd6};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd197, 8'd23, 8'd25};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd215, 8'd35, 8'd44};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd41};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd219, 8'd43, 8'd43};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd222, 8'd46, 8'd46};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd224, 8'd48, 8'd48};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd226, 8'd50, 8'd50};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd228, 8'd52, 8'd52};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd229, 8'd53, 8'd53};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd219, 8'd53, 8'd55};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd229, 8'd118, 8'd65};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd253, 8'd170, 8'd68};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd249, 8'd153, 8'd41};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd222, 8'd141, 8'd50};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd253, 8'd227, 8'd170};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd225, 8'd146, 8'd51};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd232, 8'd154, 8'd28};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd234, 8'd153, 8'd0};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd234, 8'd145, 8'd0};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd235, 8'd131, 8'd6};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd229, 8'd111, 8'd13};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd225, 8'd100, 8'd8};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd234, 8'd106, 8'd9};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd85, 8'd12};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd194, 8'd78, 8'd5};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd201, 8'd93, 8'd20};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd229, 8'd127, 8'd52};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd244, 8'd141, 8'd64};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd234, 8'd123, 8'd42};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd221, 8'd100, 8'd19};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd220, 8'd91, 8'd8};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd207, 8'd67, 8'd14};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd192, 8'd61, 8'd9};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd223, 8'd103, 8'd51};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd248, 8'd138, 8'd85};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd237, 8'd138, 8'd79};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd179, 8'd84, 8'd18};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd197, 8'd103, 8'd29};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd247, 8'd152, 8'd72};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd244, 8'd140, 8'd51};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd235, 8'd128, 8'd48};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd216, 8'd107, 8'd40};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd194, 8'd85, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd179, 8'd76, 8'd17};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd180, 8'd85, 8'd17};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd194, 8'd109, 8'd26};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd207, 8'd128, 8'd36};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd248, 8'd153, 8'd69};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd77};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd238, 8'd141, 8'd62};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd207, 8'd107, 8'd31};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd198, 8'd98, 8'd23};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd221, 8'd118, 8'd49};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd237, 8'd134, 8'd67};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd235, 8'd130, 8'd64};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd199, 8'd130, 8'd52};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd211, 8'd138, 8'd61};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd225, 8'd147, 8'd72};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd237, 8'd151, 8'd78};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd235, 8'd141, 8'd71};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd223, 8'd120, 8'd53};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd205, 8'd97, 8'd32};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd193, 8'd81, 8'd17};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd189, 8'd91, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd201, 8'd109, 8'd42};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd218, 8'd136, 8'd62};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd232, 8'd155, 8'd73};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd236, 8'd158, 8'd73};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd231, 8'd142, 8'd58};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd219, 8'd120, 8'd39};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd210, 8'd103, 8'd25};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd226, 8'd113, 8'd53};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd195, 8'd85, 8'd24};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd191, 8'd85, 8'd23};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd222, 8'd124, 8'd59};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd239, 8'd147, 8'd80};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd226, 8'd142, 8'd72};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd222, 8'd142, 8'd71};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd235, 8'd158, 8'd86};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd213, 8'd134, 8'd68};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd184, 8'd105, 8'd38};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd170, 8'd87, 8'd17};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd188, 8'd104, 8'd31};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd220, 8'd133, 8'd54};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd234, 8'd143, 8'd62};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd225, 8'd133, 8'd48};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd215, 8'd121, 8'd34};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd194, 8'd88, 8'd26};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd191, 8'd97, 8'd33};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd198, 8'd114, 8'd50};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd232, 8'd144, 8'd81};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd229, 8'd129, 8'd67};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd219, 8'd112, 8'd42};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd201, 8'd99, 8'd15};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd208, 8'd113, 8'd19};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd211, 8'd131, 8'd10};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd240, 8'd148, 8'd3};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd229, 8'd131, 8'd0};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd200, 8'd122, 8'd11};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd222, 8'd179, 8'd136};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd245, 8'd223, 8'd199};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd232, 8'd152, 8'd67};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd227, 8'd145, 8'd20};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd255, 8'd171, 8'd56};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd253, 8'd127, 8'd77};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd203, 8'd50, 8'd45};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd231, 8'd63, 8'd52};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd225, 8'd45, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd235, 8'd47, 8'd48};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd222, 8'd44, 8'd44};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd221, 8'd43, 8'd43};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd215, 8'd39, 8'd39};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd209, 8'd33, 8'd33};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd200, 8'd26, 8'd25};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd190, 8'd16, 8'd15};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd181, 8'd9, 8'd7};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd176, 8'd4, 8'd2};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd158, 8'd4, 8'd4};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd161, 8'd0, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd169, 8'd1, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd156, 8'd0, 8'd0};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd148, 8'd4, 8'd4};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd170, 8'd45, 8'd13};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd247, 8'd133, 8'd47};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd250, 8'd139, 8'd8};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd249, 8'd127, 8'd16};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd209, 8'd130, 8'd53};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd205, 8'd175, 8'd141};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd128: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd234, 8'd218, 8'd202};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd201, 8'd127, 8'd42};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd244, 8'd135, 8'd34};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd235, 8'd151, 8'd27};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd248, 8'd149, 8'd32};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd230, 8'd81, 8'd51};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd146, 8'd4, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd164, 8'd10, 8'd8};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd161, 8'd7, 8'd5};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd160, 8'd2, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd161, 8'd0, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd166, 8'd1, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd175, 8'd6, 8'd3};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd186, 8'd12, 8'd11};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd191, 8'd17, 8'd16};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd206, 8'd32, 8'd41};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd219, 8'd46, 8'd42};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd216, 8'd40, 8'd27};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd224, 8'd46, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd221, 8'd41, 8'd42};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd216, 8'd39, 8'd45};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd229, 8'd57, 8'd55};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd216, 8'd48, 8'd37};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd216, 8'd83, 8'd52};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd255, 8'd165, 8'd75};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd238, 8'd159, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd225, 8'd138, 8'd32};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd248, 8'd190, 8'd142};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd252, 8'd226, 8'd167};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd216, 8'd158, 8'd61};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd249, 8'd146, 8'd0};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd242, 8'd140, 8'd0};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd234, 8'd133, 8'd1};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd230, 8'd127, 8'd9};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd229, 8'd120, 8'd19};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd229, 8'd109, 8'd22};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd224, 8'd94, 8'd16};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd220, 8'd84, 8'd10};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd201, 8'd88, 8'd18};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd159, 8'd48, 8'd0};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd181, 8'd81, 8'd22};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd248, 8'd169, 8'd74};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd254, 8'd191, 8'd50};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd251, 8'd177, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd210, 8'd102, 8'd0};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd217, 8'd77, 8'd16};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd177, 8'd50, 8'd7};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd142, 8'd57, 8'd0};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd239, 8'd190, 8'd114};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd138};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd249, 8'd166, 8'd112};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd140, 8'd39, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd242, 8'd160, 8'd78};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd243, 8'd190, 8'd78};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd228, 8'd201, 8'd96};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd206, 8'd96, 8'd21};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd208, 8'd86, 8'd21};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd142, 8'd56, 8'd0};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd177, 8'd89, 8'd17};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd238, 8'd166, 8'd84};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd242, 8'd198, 8'd101};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd251, 8'd199, 8'd100};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd248, 8'd195, 8'd91};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd253, 8'd202, 8'd110};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd124};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd211, 8'd149, 8'd66};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd186, 8'd114, 8'd16};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd249, 8'd180, 8'd63};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd253, 8'd200, 8'd72};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd235, 8'd197, 8'd64};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd64};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd249, 8'd192, 8'd87};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd249, 8'd209, 8'd113};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd249, 8'd215, 8'd107};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd243, 8'd194, 8'd101};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd243, 8'd175, 8'd114};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd133, 8'd58, 8'd1};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd179, 8'd111, 8'd28};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd224, 8'd159, 8'd69};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd247, 8'd179, 8'd82};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd93};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd252, 8'd200, 8'd99};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd240, 8'd200, 8'd105};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd232, 8'd193, 8'd98};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd242, 8'd190, 8'd88};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd212, 8'd146, 8'd34};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd194, 8'd105, 8'd45};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd175, 8'd69, 8'd7};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd209, 8'd115, 8'd41};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd241, 8'd186, 8'd95};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd242, 8'd202, 8'd107};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd122};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd142};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd233, 8'd219, 8'd148};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd227, 8'd205, 8'd155};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd239, 8'd194, 8'd139};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd193, 8'd124, 8'd57};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd182, 8'd110, 8'd26};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd241, 8'd183, 8'd84};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd104};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd255, 8'd197, 8'd105};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd195, 8'd102, 8'd22};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd181, 8'd104, 8'd50};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd163, 8'd92, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd243, 8'd177, 8'd103};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd254, 8'd189, 8'd105};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd246, 8'd173, 8'd81};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd204, 8'd113, 8'd22};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd212, 8'd102, 8'd15};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd209, 8'd87, 8'd4};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd216, 8'd120, 8'd17};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd217, 8'd123, 8'd9};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd216, 8'd125, 8'd0};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd233, 8'd142, 8'd1};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd223, 8'd144, 8'd15};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd226, 8'd174, 8'd88};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd253, 8'd242, 8'd210};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd227, 8'd189, 8'd118};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd216, 8'd141, 8'd48};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd243, 8'd146, 8'd31};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd57};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd209, 8'd76, 8'd31};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd217, 8'd42, 8'd47};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd228, 8'd48, 8'd57};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd220, 8'd66, 8'd54};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd225, 8'd53, 8'd51};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd218, 8'd44, 8'd43};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd207, 8'd31, 8'd31};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd195, 8'd16, 8'd19};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd183, 8'd7, 8'd10};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd176, 8'd3, 8'd5};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd172, 8'd3, 8'd6};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd170, 8'd6, 8'd7};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd153, 8'd7, 8'd0};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd147, 8'd0, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd163, 8'd9, 8'd7};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd163, 8'd8, 8'd14};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd167, 8'd15, 8'd12};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd172, 8'd30, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd241, 8'd113, 8'd24};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd150, 8'd21};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd240, 8'd133, 8'd17};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd218, 8'd134, 8'd48};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd193, 8'd146, 8'd100};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd129: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd225, 8'd211, 8'd200};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd190, 8'd120, 8'd34};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd246, 8'd141, 8'd36};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd26};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd234, 8'd139, 8'd23};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd204, 8'd58, 8'd35};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd145, 8'd3, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd163, 8'd5, 8'd4};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd161, 8'd1, 8'd1};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd159, 8'd0, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd161, 8'd0, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd165, 8'd0, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd174, 8'd6, 8'd3};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd183, 8'd14, 8'd11};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd190, 8'd18, 8'd16};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd202, 8'd28, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd216, 8'd43, 8'd39};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd217, 8'd41, 8'd28};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd41};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd226, 8'd46, 8'd49};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd220, 8'd43, 8'd49};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd231, 8'd59, 8'd57};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd221, 8'd55, 8'd41};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd227, 8'd98, 8'd56};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd67};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd26};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd229, 8'd147, 8'd47};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd254, 8'd203, 8'd156};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd253, 8'd231, 8'd194};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd234, 8'd186, 8'd101};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd217, 8'd147, 8'd23};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd248, 8'd146, 8'd2};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd239, 8'd137, 8'd1};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd228, 8'd126, 8'd2};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd222, 8'd118, 8'd7};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd222, 8'd112, 8'd14};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd226, 8'd106, 8'd19};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd228, 8'd99, 8'd18};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd226, 8'd93, 8'd16};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd210, 8'd87, 8'd20};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd173, 8'd56, 8'd3};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd150, 8'd51, 8'd0};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd233, 8'd163, 8'd77};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd244, 8'd193, 8'd66};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd68};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd200, 8'd102, 8'd11};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd203, 8'd73, 8'd24};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd157, 8'd38, 8'd16};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd172, 8'd93, 8'd50};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd151};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd152};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd220, 8'd142, 8'd96};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd122, 8'd28, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd230, 8'd158, 8'd76};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd242, 8'd200, 8'd88};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd117};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd192, 8'd82, 8'd5};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd182, 8'd68, 8'd0};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd170, 8'd96, 8'd11};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd231, 8'd155, 8'd69};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd255, 8'd185, 8'd89};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd91};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd238, 8'd171, 8'd58};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd237, 8'd164, 8'd59};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd238, 8'd167, 8'd75};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd244, 8'd171, 8'd92};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd218, 8'd136, 8'd60};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd200, 8'd110, 8'd24};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd239, 8'd153, 8'd54};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd227, 8'd158, 8'd54};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd223, 8'd170, 8'd66};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd68};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd204, 8'd101};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd231, 8'd177, 8'd81};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd220, 8'd166, 8'd58};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd247, 8'd178, 8'd83};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd205, 8'd124, 8'd59};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd155, 8'd76, 8'd10};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd235, 8'd169, 8'd75};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd87};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd249, 8'd186, 8'd70};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd237, 8'd167, 8'd53};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd222, 8'd157, 8'd53};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd212, 8'd157, 8'd66};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd246, 8'd199, 8'd111};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd113};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd243, 8'd181, 8'd80};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd199, 8'd118, 8'd55};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd176, 8'd79, 8'd11};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd212, 8'd128, 8'd42};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd246, 8'd202, 8'd97};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd247, 8'd213, 8'd115};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd255, 8'd213, 8'd141};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd178};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd202};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd190};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd171};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd236, 8'd173, 8'd119};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd193, 8'd128, 8'd60};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd217, 8'd162, 8'd79};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd247, 8'd198, 8'd105};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd106};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd211, 8'd136, 8'd45};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd140, 8'd65, 8'd0};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd177, 8'd108, 8'd33};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd111};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd255, 8'd193, 8'd102};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd223, 8'd147, 8'd53};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd198, 8'd104, 8'd14};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd207, 8'd95, 8'd11};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd218, 8'd93, 8'd13};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd214, 8'd111, 8'd10};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd220, 8'd122, 8'd13};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd228, 8'd136, 8'd13};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd223, 8'd132, 8'd0};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd210, 8'd128, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd206, 8'd146, 8'd48};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd228, 8'd198, 8'd146};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd238, 8'd208, 8'd146};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd220, 8'd150, 8'd62};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd244, 8'd148, 8'd35};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd58};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd222, 8'd92, 8'd42};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd217, 8'd45, 8'd43};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd227, 8'd46, 8'd51};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd220, 8'd60, 8'd46};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd216, 8'd44, 8'd42};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd210, 8'd36, 8'd35};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd200, 8'd24, 8'd24};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd191, 8'd12, 8'd15};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd180, 8'd4, 8'd7};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd174, 8'd1, 8'd3};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd171, 8'd2, 8'd5};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd168, 8'd4, 8'd5};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd180, 8'd6, 8'd8};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd165, 8'd0, 8'd0};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd168, 8'd0, 8'd3};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd167, 8'd0, 8'd12};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd166, 8'd10, 8'd14};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd162, 8'd32, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd222, 8'd118, 8'd29};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd245, 8'd160, 8'd31};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd246, 8'd143, 8'd15};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd226, 8'd143, 8'd51};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd203, 8'd155, 8'd109};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd130: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd238, 8'd221, 8'd211};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd191, 8'd122, 8'd31};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd245, 8'd144, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd231, 8'd153, 8'd19};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd238, 8'd141, 8'd24};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd197, 8'd47, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd162, 8'd14, 8'd14};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd166, 8'd0, 8'd2};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd164, 8'd0, 8'd0};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd162, 8'd0, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd162, 8'd0, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd165, 8'd0, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd171, 8'd6, 8'd2};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd178, 8'd13, 8'd9};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd182, 8'd17, 8'd13};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd195, 8'd20, 8'd27};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd210, 8'd35, 8'd32};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd216, 8'd39, 8'd29};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd227, 8'd48, 8'd41};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd228, 8'd49, 8'd52};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd222, 8'd48, 8'd50};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd229, 8'd60, 8'd53};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd230, 8'd65, 8'd46};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd243, 8'd123, 8'd60};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd250, 8'd156, 8'd56};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd224, 8'd145, 8'd26};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd233, 8'd164, 8'd71};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd184};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd217};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd241, 8'd178, 8'd109};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd221, 8'd140, 8'd22};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd234, 8'd148, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd245, 8'd142, 8'd14};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd233, 8'd130, 8'd9};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd220, 8'd116, 8'd3};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd213, 8'd105, 8'd4};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd216, 8'd103, 8'd9};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd223, 8'd103, 8'd16};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd229, 8'd103, 8'd19};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd232, 8'd101, 8'd19};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd227, 8'd87, 8'd26};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd189, 8'd63, 8'd13};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd127, 8'd31, 8'd0};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd189, 8'd131, 8'd57};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd244, 8'd211, 8'd108};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd117};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd202, 8'd121, 8'd55};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd178, 8'd63, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd132, 8'd31, 8'd23};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd214, 8'd149, 8'd121};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd189};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd171};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd189, 8'd114, 8'd82};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd114, 8'd29, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd222, 8'd163, 8'd93};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd243, 8'd219, 8'd119};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd216, 8'd125};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd162, 8'd57, 8'd0};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd149, 8'd52, 8'd0};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd207, 8'd157, 8'd70};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd253, 8'd199, 8'd103};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd244, 8'd181, 8'd75};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd236, 8'd174, 8'd53};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd224, 8'd135, 8'd15};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd212, 8'd114, 8'd5};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd208, 8'd113, 8'd19};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd211, 8'd118, 8'd40};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd203, 8'd102, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd194, 8'd86, 8'd14};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd199, 8'd97, 8'd23};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd166, 8'd82, 8'd12};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd182, 8'd113, 8'd48};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd251, 8'd194, 8'd78};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd252, 8'd193, 8'd103};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd219, 8'd156, 8'd76};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd185, 8'd112, 8'd18};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd190, 8'd104, 8'd19};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd163, 8'd73, 8'd13};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd215, 8'd141, 8'd76};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd243, 8'd190, 8'd94};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd245, 8'd206, 8'd75};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd228, 8'd171, 8'd42};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd211, 8'd132, 8'd14};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd194, 8'd108, 8'd9};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd162, 8'd85, 8'd3};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd210, 8'd147, 8'd70};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd246, 8'd191, 8'd108};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd254, 8'd201, 8'd109};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd228, 8'd155, 8'd87};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd178, 8'd92, 8'd19};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd211, 8'd140, 8'd52};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd254, 8'd221, 8'd118};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd241, 8'd218, 8'd125};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd223, 8'd179, 8'd118};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd216, 8'd171, 8'd140};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd223, 8'd198, 8'd178};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd190};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd184};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd255, 8'd210, 8'd167};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd194, 8'd131, 8'd80};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd173, 8'd118, 8'd53};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd224, 8'd173, 8'd90};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd251, 8'd198, 8'd102};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd225, 8'd166, 8'd62};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd139, 8'd72, 8'd0};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd213, 8'd148, 8'd58};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd110};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd253, 8'd181, 8'd83};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd202, 8'd119, 8'd23};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd202, 8'd102, 8'd14};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd209, 8'd94, 8'd13};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd222, 8'd99, 8'd22};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd216, 8'd99, 8'd3};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd214, 8'd108, 8'd6};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd224, 8'd130, 8'd17};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd214, 8'd126, 8'd0};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd218, 8'd133, 8'd4};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd212, 8'd136, 8'd24};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd203, 8'd147, 8'd62};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd155};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd253, 8'd235, 8'd187};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd226, 8'd163, 8'd86};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd244, 8'd149, 8'd41};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd255, 8'd159, 8'd53};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd237, 8'd113, 8'd53};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd214, 8'd48, 8'd36};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd223, 8'd41, 8'd40};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd217, 8'd47, 8'd32};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd203, 8'd31, 8'd29};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd198, 8'd24, 8'd23};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd191, 8'd15, 8'd15};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd184, 8'd5, 8'd8};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd176, 8'd0, 8'd3};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd172, 8'd0, 8'd1};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd169, 8'd0, 8'd3};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd167, 8'd3, 8'd4};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd173, 8'd2, 8'd8};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd175, 8'd0, 8'd6};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd189, 8'd4, 8'd18};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd194, 8'd8, 8'd29};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd178, 8'd7, 8'd16};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd162, 8'd18, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd214, 8'd102, 8'd28};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd250, 8'd160, 8'd46};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd237, 8'd143, 8'd7};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd221, 8'd145, 8'd47};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd207, 8'd160, 8'd114};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd131: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd246, 8'd223, 8'd209};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd192, 8'd116, 8'd18};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd244, 8'd138, 8'd16};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd233, 8'd152, 8'd9};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd247, 8'd144, 8'd23};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd190, 8'd31, 8'd12};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd164, 8'd6, 8'd7};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd174, 8'd4, 8'd7};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd172, 8'd2, 8'd5};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd168, 8'd0, 8'd0};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd166, 8'd0, 8'd0};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd165, 8'd0, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd167, 8'd4, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd170, 8'd7, 8'd2};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd172, 8'd10, 8'd5};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd185, 8'd8, 8'd14};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd201, 8'd23, 8'd21};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd210, 8'd32, 8'd22};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd220, 8'd41, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd225, 8'd46, 8'd49};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd218, 8'd44, 8'd46};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd221, 8'd55, 8'd43};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd233, 8'd74, 8'd45};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd255, 8'd147, 8'd62};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd243, 8'd150, 8'd46};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd218, 8'd142, 8'd32};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd240, 8'd185, 8'd103};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd251, 8'd240, 8'd234};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd247, 8'd191, 8'd134};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd233, 8'd141, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd234, 8'd128, 8'd0};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd248, 8'd143, 8'd0};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd234, 8'd133, 8'd19};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd225, 8'd123, 8'd13};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd216, 8'd110, 8'd8};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd211, 8'd102, 8'd7};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd216, 8'd102, 8'd13};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd224, 8'd104, 8'd17};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd229, 8'd105, 8'd19};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd230, 8'd104, 8'd17};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd242, 8'd92, 8'd33};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd202, 8'd70, 8'd21};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd138, 8'd41, 8'd0};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd134, 8'd80, 8'd20};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd253, 8'd228, 8'd148};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd151};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd225, 8'd162, 8'd111};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd154, 8'd60, 8'd35};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd127, 8'd47, 8'd24};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd247, 8'd198, 8'd158};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd255, 8'd241, 8'd191};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd249, 8'd207, 8'd167};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd180, 8'd105, 8'd84};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd136, 8'd55, 8'd36};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd234, 8'd185, 8'd142};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd250, 8'd240, 8'd169};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd165};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd154, 8'd60, 8'd22};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd148, 8'd75, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd246, 8'd227, 8'd158};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd254, 8'd227, 8'd146};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd243, 8'd196, 8'd104};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd218, 8'd154, 8'd48};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd229, 8'd128, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd237, 8'd129, 8'd18};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd232, 8'd130, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd229, 8'd128, 8'd46};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd225, 8'd118, 8'd46};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd221, 8'd109, 8'd45};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd209, 8'd104, 8'd47};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd161, 8'd74, 8'd31};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd187, 8'd113, 8'd84};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd247, 8'd220, 8'd133};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd247, 8'd211, 8'd151};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd232, 8'd181, 8'd128};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd190, 8'd121, 8'd54};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd173, 8'd91, 8'd31};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd162, 8'd87, 8'd47};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd254, 8'd206, 8'd157};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd243, 8'd225, 8'd143};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd242, 8'd212, 8'd102};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd226, 8'd169, 8'd62};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd223, 8'd133, 8'd37};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd221, 8'd115, 8'd37};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd176, 8'd78, 8'd13};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd179, 8'd104, 8'd37};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd241, 8'd186, 8'd104};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd253, 8'd207, 8'd113};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd246, 8'd183, 8'd106};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd166, 8'd87, 8'd20};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd197, 8'd134, 8'd67};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd160};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd238, 8'd219, 8'd151};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd183, 8'd142, 8'd88};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd152, 8'd106, 8'd57};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd168, 8'd143, 8'd87};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd243, 8'd215, 8'd152};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd161};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd158};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd201, 8'd130, 8'd84};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd159, 8'd90, 8'd31};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd204, 8'd143, 8'd63};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd247, 8'd194, 8'd90};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd239, 8'd188, 8'd71};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd197, 8'd139, 8'd39};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd252, 8'd193, 8'd91};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd92};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd223, 8'd148, 8'd46};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd198, 8'd110, 8'd13};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd212, 8'd111, 8'd21};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd218, 8'd103, 8'd23};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd224, 8'd102, 8'd27};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd225, 8'd100, 8'd7};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd210, 8'd100, 8'd3};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd206, 8'd113, 8'd9};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd208, 8'd122, 8'd3};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd223, 8'd136, 8'd5};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd222, 8'd134, 8'd8};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd207, 8'd130, 8'd16};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd230, 8'd160, 8'd62};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd243, 8'd224, 8'd192};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd231, 8'd173, 8'd109};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd237, 8'd144, 8'd40};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd252, 8'd154, 8'd43};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd248, 8'd131, 8'd61};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd208, 8'd49, 8'd27};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd216, 8'd33, 8'd29};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd208, 8'd30, 8'd16};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd191, 8'd19, 8'd17};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd189, 8'd15, 8'd14};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd184, 8'd8, 8'd8};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd181, 8'd2, 8'd5};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd175, 8'd0, 8'd2};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd172, 8'd0, 8'd1};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd170, 8'd1, 8'd4};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd168, 8'd4, 8'd5};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd155, 8'd12, 8'd4};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd165, 8'd10, 8'd5};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd182, 8'd9, 8'd11};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd203, 8'd17, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd197, 8'd11, 8'd22};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd185, 8'd15, 8'd2};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd226, 8'd81, 8'd26};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd136, 8'd49};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd224, 8'd146, 8'd12};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd214, 8'd149, 8'd55};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd208, 8'd166, 8'd124};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd132: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd246, 8'd215, 8'd194};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd193, 8'd114, 8'd13};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd148, 8'd27};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd252, 8'd166, 8'd27};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd252, 8'd143, 8'd22};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd182, 8'd16, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd172, 8'd5, 8'd0};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd183, 8'd10, 8'd14};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd181, 8'd8, 8'd12};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd175, 8'd5, 8'd6};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd171, 8'd3, 8'd3};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd168, 8'd0, 8'd0};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd166, 8'd1, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd165, 8'd2, 8'd0};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd165, 8'd2, 8'd0};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd178, 8'd0, 8'd3};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd191, 8'd12, 8'd8};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd202, 8'd21, 8'd14};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd210, 8'd28, 8'd25};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd216, 8'd37, 8'd41};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd209, 8'd37, 8'd37};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd209, 8'd46, 8'd27};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd236, 8'd79, 8'd44};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd58};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd239, 8'd144, 8'd38};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd219, 8'd143, 8'd47};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd247, 8'd208, 8'd141};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd226, 8'd214, 8'd174};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd212, 8'd157, 8'd56};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd240, 8'd144, 8'd5};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd255, 8'd149, 8'd13};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd245, 8'd132, 8'd14};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd224, 8'd127, 8'd20};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd220, 8'd118, 8'd17};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd216, 8'd109, 8'd13};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd216, 8'd105, 8'd15};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd221, 8'd105, 8'd18};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd226, 8'd106, 8'd19};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd226, 8'd105, 8'd16};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd224, 8'd103, 8'd12};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd244, 8'd96, 8'd32};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd219, 8'd86, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd162, 8'd62, 8'd13};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd109, 8'd49, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd237, 8'd208, 8'd148};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd170};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd249, 8'd197, 8'd147};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd146, 8'd71, 8'd32};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd147, 8'd85, 8'd26};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd151};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd253, 8'd229, 8'd155};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd235, 8'd189, 8'd139};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd191, 8'd112, 8'd95};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd171, 8'd88, 8'd82};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd253, 8'd208, 8'd187};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd255, 8'd253, 8'd210};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd215};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd148, 8'd68, 8'd57};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd169, 8'd116, 8'd98};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd249, 8'd251, 8'd211};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd196};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd245, 8'd211, 8'd147};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd210, 8'd151, 8'd71};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd230, 8'd129, 8'd49};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd238, 8'd136, 8'd26};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd238, 8'd140, 8'd41};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd229, 8'd135, 8'd48};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd221, 8'd124, 8'd47};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd225, 8'd122, 8'd55};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd217, 8'd120, 8'd69};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd165, 8'd86, 8'd55};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd190, 8'd127, 8'd112};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd246, 8'd251, 8'd195};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd219};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd236, 8'd208, 8'd184};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd212, 8'd164, 8'd124};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd213, 8'd153, 8'd117};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd183, 8'd131, 8'd117};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd229, 8'd211, 8'd187};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd252, 8'd255, 8'd211};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd161};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd232, 8'd171, 8'd104};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd240, 8'd142, 8'd79};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd255, 8'd140, 8'd86};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd215, 8'd108, 8'd56};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd164, 8'd83, 8'd20};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd247, 8'd191, 8'd104};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd239, 8'd196, 8'd91};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd240, 8'd179, 8'd98};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd152, 8'd76, 8'd18};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd189, 8'd127, 8'd90};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd199};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd254, 8'd235, 8'd195};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd212, 8'd169, 8'd114};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd179, 8'd131, 8'd46};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd198, 8'd168, 8'd54};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd249, 8'd202, 8'd122};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd247, 8'd193, 8'd121};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd239, 8'd171, 8'd110};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd227, 8'd146, 8'd90};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd191, 8'd103, 8'd40};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd189, 8'd108, 8'd29};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd230, 8'd166, 8'd66};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd254, 8'd205, 8'd87};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd242, 8'd197, 8'd96};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd107};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd239, 8'd174, 8'd74};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd201, 8'd123, 8'd23};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd211, 8'd118, 8'd23};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd220, 8'd116, 8'd27};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd225, 8'd114, 8'd32};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd224, 8'd108, 8'd31};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd235, 8'd110, 8'd18};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd216, 8'd105, 8'd13};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd195, 8'd103, 8'd2};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd205, 8'd120, 8'd3};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd211, 8'd123, 8'd0};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd219, 8'd129, 8'd0};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd232, 8'd149, 8'd19};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd213, 8'd137, 8'd17};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd214, 8'd192, 8'd153};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd235, 8'd182, 8'd128};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd231, 8'd135, 8'd33};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd246, 8'd149, 8'd32};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd248, 8'd142, 8'd58};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd203, 8'd56, 8'd23};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd206, 8'd27, 8'd20};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd201, 8'd19, 8'd8};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd188, 8'd16, 8'd14};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd187, 8'd13, 8'd12};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd184, 8'd8, 8'd8};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd183, 8'd4, 8'd7};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd179, 8'd3, 8'd6};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd176, 8'd3, 8'd5};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd174, 8'd5, 8'd8};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd171, 8'd7, 8'd8};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd167, 8'd15, 8'd2};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd186, 8'd28, 8'd16};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd191, 8'd23, 8'd14};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd191, 8'd17, 8'd18};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd163, 8'd0, 8'd0};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd151, 8'd0, 8'd0};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd201, 8'd70, 8'd28};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd255, 8'd141, 8'd71};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd231, 8'd174, 8'd67};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd225, 8'd177, 8'd103};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd226, 8'd193, 8'd162};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd133: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd232, 8'd207, 8'd185};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd185, 8'd111, 8'd22};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd248, 8'd145, 8'd44};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd240, 8'd161, 8'd42};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd225, 8'd124, 8'd16};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd168, 8'd9, 8'd0};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd182, 8'd21, 8'd11};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd184, 8'd14, 8'd17};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd182, 8'd12, 8'd15};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd180, 8'd10, 8'd11};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd177, 8'd7, 8'd8};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd174, 8'd4, 8'd4};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd171, 8'd2, 8'd0};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd170, 8'd1, 8'd0};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd169, 8'd0, 8'd0};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd178, 8'd0, 8'd1};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd188, 8'd6, 8'd3};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd196, 8'd14, 8'd10};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd199, 8'd17, 8'd16};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd207, 8'd28, 8'd32};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd198, 8'd29, 8'd26};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd200, 8'd40, 8'd16};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd241, 8'd88, 8'd46};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd254, 8'd168, 8'd49};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd236, 8'd140, 8'd37};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd227, 8'd152, 8'd71};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd253, 8'd228, 8'd174};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd227, 8'd211, 8'd159};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd196, 8'd155, 8'd41};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd228, 8'd157, 8'd13};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd41};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd248, 8'd143, 8'd38};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd224, 8'd129, 8'd21};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd220, 8'd121, 8'd19};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd218, 8'd111, 8'd15};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd220, 8'd106, 8'd17};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd225, 8'd107, 8'd20};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd228, 8'd108, 8'd21};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd225, 8'd107, 8'd17};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd222, 8'd105, 8'd12};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd232, 8'd99, 8'd22};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd229, 8'd102, 8'd35};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd182, 8'd75, 8'd19};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd125, 8'd49, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd196, 8'd149, 8'd97};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd164};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd142};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd160, 8'd97, 8'd28};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd183, 8'd127, 8'd40};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd255, 8'd221, 8'd124};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd240, 8'd210, 8'd114};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd220, 8'd163, 8'd96};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd206, 8'd115, 8'd84};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd188, 8'd96, 8'd83};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd185};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd252, 8'd251, 8'd207};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd215};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd149, 8'd74, 8'd69};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd199, 8'd149, 8'd142};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd240, 8'd246, 8'd218};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd215};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd234, 8'd202, 8'd153};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd216, 8'd161, 8'd97};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd239, 8'd140, 8'd75};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd243, 8'd146, 8'd49};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd239, 8'd150, 8'd58};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd233, 8'd147, 8'd62};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd229, 8'd138, 8'd59};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd236, 8'd142, 8'd68};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd236, 8'd145, 8'd88};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd188, 8'd113, 8'd81};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd208, 8'd149, 8'd135};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd248, 8'd255, 8'd216};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd254, 8'd255, 8'd235};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd252, 8'd236, 8'd220};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd235, 8'd201, 8'd166};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd217, 8'd170, 8'd142};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd202, 8'd161, 8'd157};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd238, 8'd228, 8'd219};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd243, 8'd255, 8'd225};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd175};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd220, 8'd158, 8'd107};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd243, 8'd147, 8'd97};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd254, 8'd142, 8'd96};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd207, 8'd102, 8'd54};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd140, 8'd61, 8'd0};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd242, 8'd185, 8'd95};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd239, 8'd193, 8'd82};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd241, 8'd176, 8'd96};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd160, 8'd80, 8'd27};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd201, 8'd138, 8'd107};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd209};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd210};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd146};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd239, 8'd180, 8'd76};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd80};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd108};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd236, 8'd177, 8'd87};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd208, 8'd140, 8'd59};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd243, 8'd156, 8'd85};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd223, 8'd124, 8'd57};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd171, 8'd77, 8'd5};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd186, 8'd116, 8'd31};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd209, 8'd115};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd247, 8'd211, 8'd125};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd247, 8'd201, 8'd115};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd219, 8'd158, 8'd69};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd205, 8'd125, 8'd36};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd222, 8'd128, 8'd38};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd220, 8'd119, 8'd31};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd225, 8'd121, 8'd34};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd225, 8'd119, 8'd33};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd237, 8'd118, 8'd26};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd213, 8'd109, 8'd14};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd192, 8'd100, 8'd0};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd213, 8'd128, 8'd9};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd223, 8'd137, 8'd2};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd232, 8'd149, 8'd11};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd242, 8'd169, 8'd38};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd193, 8'd131, 8'd10};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd208, 8'd191, 8'd148};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd246, 8'd192, 8'd145};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd228, 8'd129, 8'd28};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd243, 8'd147, 8'd24};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd245, 8'd148, 8'd54};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd202, 8'd69, 8'd28};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd202, 8'd31, 8'd23};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd200, 8'd17, 8'd13};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd192, 8'd20, 8'd18};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd192, 8'd18, 8'd17};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd191, 8'd15, 8'd15};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd191, 8'd12, 8'd15};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd187, 8'd11, 8'd14};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd184, 8'd11, 8'd13};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd180, 8'd11, 8'd14};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd177, 8'd13, 8'd14};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd191, 8'd3, 8'd4};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd195, 8'd16, 8'd12};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd165, 8'd4, 8'd0};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd161, 8'd22, 8'd17};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd154, 8'd40, 8'd40};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd167, 8'd80, 8'd71};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd203, 8'd140, 8'd107};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd238, 8'd191, 8'd139};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd159};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd250, 8'd221, 8'd181};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd249, 8'd230, 8'd216};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd134: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd218, 8'd215, 8'd200};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd196, 8'd141, 8'd74};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd236, 8'd152, 8'd82};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd218, 8'd158, 8'd72};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd202, 8'd120, 8'd36};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd160, 8'd19, 8'd12};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd167, 8'd26, 8'd19};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd176, 8'd12, 8'd13};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd176, 8'd12, 8'd13};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd177, 8'd11, 8'd11};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd180, 8'd10, 8'd11};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd182, 8'd10, 8'd10};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd182, 8'd8, 8'd7};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd182, 8'd6, 8'd6};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd182, 8'd6, 8'd6};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd186, 8'd3, 8'd7};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd191, 8'd7, 8'd5};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd196, 8'd13, 8'd9};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd193, 8'd10, 8'd12};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd201, 8'd22, 8'd28};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd194, 8'd25, 8'd20};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd195, 8'd37, 8'd10};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd249, 8'd98, 8'd51};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd244, 8'd165, 8'd38};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd235, 8'd137, 8'd38};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd237, 8'd162, 8'd95};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd201};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd251, 8'd231, 8'd194};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd214, 8'd193, 8'd104};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd213, 8'd177, 8'd54};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd239, 8'd175, 8'd49};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd250, 8'd163, 8'd47};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd231, 8'd141, 8'd27};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd225, 8'd128, 8'd21};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd219, 8'd113, 8'd13};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd217, 8'd104, 8'd12};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd221, 8'd103, 8'd15};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd225, 8'd107, 8'd19};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd225, 8'd110, 8'd19};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd224, 8'd111, 8'd17};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd218, 8'd103, 8'd14};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd222, 8'd103, 8'd23};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd199, 8'd85, 8'd22};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd154, 8'd58, 8'd7};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd158, 8'd88, 8'd37};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd249, 8'd198, 8'd133};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd254, 8'd204, 8'd117};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd181, 8'd128, 8'd24};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd215, 8'd159, 8'd66};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd248, 8'd207, 8'd102};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd237, 8'd196, 8'd90};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd205, 8'd137, 8'd52};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd210, 8'd106, 8'd55};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd172, 8'd73, 8'd34};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd234, 8'd185, 8'd129};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd235, 8'd236, 8'd160};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd176};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd168, 8'd87, 8'd58};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd199, 8'd139, 8'd115};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd211};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd205};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd248, 8'd207, 8'd153};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd232, 8'd172, 8'd102};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd254, 8'd153, 8'd83};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd240, 8'd143, 8'd62};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd227, 8'd138, 8'd58};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd226, 8'd139, 8'd60};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd231, 8'd140, 8'd59};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd234, 8'd137, 8'd58};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd227, 8'd133, 8'd69};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd178, 8'd99, 8'd60};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd195, 8'd130, 8'd110};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd255, 8'd248, 8'd193};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd212};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd208};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd244, 8'd204, 8'd153};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd206, 8'd153, 8'd111};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd201, 8'd149, 8'd135};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd228};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd246, 8'd243, 8'd202};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd157};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd206, 8'd149, 8'd80};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd244, 8'd157, 8'd90};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd235, 8'd135, 8'd75};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd179, 8'd86, 8'd29};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd155, 8'd80, 8'd13};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd250, 8'd190, 8'd102};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd104};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd248, 8'd174, 8'd103};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd160, 8'd78, 8'd20};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd205, 8'd144, 8'd90};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd255, 8'd237, 8'd179};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd253, 8'd232, 8'd167};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd233, 8'd177, 8'd103};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd218, 8'd142, 8'd54};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd89};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd104};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd236, 8'd182, 8'd84};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd205, 8'd146, 8'd52};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd231, 8'd153, 8'd70};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd234, 8'd137, 8'd68};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd181, 8'd86, 8'd28};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd155, 8'd90, 8'd34};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd159};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd249, 8'd222, 8'd155};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd138};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd214, 8'd154, 8'd81};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd224, 8'd145, 8'd66};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd225, 8'd133, 8'd48};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd228, 8'd128, 8'd40};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd225, 8'd126, 8'd33};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd223, 8'd126, 8'd32};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd227, 8'd118, 8'd23};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd210, 8'd112, 8'd13};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd203, 8'd115, 8'd7};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd226, 8'd141, 8'd16};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd244, 8'd161, 8'd23};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd242, 8'd169, 8'd31};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd225, 8'd171, 8'd47};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd198, 8'd162, 8'd52};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd234, 8'd222, 8'd180};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd160};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd231, 8'd128, 8'd27};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd246, 8'd151, 8'd21};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd242, 8'd153, 8'd51};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd208, 8'd86, 8'd39};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd203, 8'd38, 8'd32};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd203, 8'd23, 8'd26};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd200, 8'd28, 8'd26};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd200, 8'd26, 8'd25};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd200, 8'd24, 8'd24};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd201, 8'd22, 8'd25};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd196, 8'd20, 8'd23};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd192, 8'd19, 8'd21};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd187, 8'd18, 8'd21};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd183, 8'd19, 8'd20};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd182, 8'd1, 8'd16};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd185, 8'd26, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd152, 8'd30, 8'd25};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd179, 8'd98, 8'd95};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd221, 8'd172, 8'd176};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd135: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd255, 8'd217, 8'd168};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd162};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd246, 8'd202, 8'd141};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd233, 8'd168, 8'd104};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd185, 8'd60, 8'd64};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd159, 8'd35, 8'd33};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd167, 8'd7, 8'd7};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd171, 8'd8, 8'd9};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd175, 8'd11, 8'd10};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd181, 8'd13, 8'd13};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd187, 8'd13, 8'd14};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd192, 8'd14, 8'd14};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd193, 8'd13, 8'd14};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd196, 8'd13, 8'd15};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd193, 8'd9, 8'd11};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd194, 8'd10, 8'd8};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd198, 8'd15, 8'd11};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd191, 8'd8, 8'd10};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd198, 8'd21, 8'd27};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd193, 8'd24, 8'd19};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd195, 8'd37, 8'd8};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd105, 8'd54};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd235, 8'd161, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd235, 8'd136, 8'd42};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd245, 8'd169, 8'd111};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd251, 8'd215};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd252, 8'd242, 8'd183};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd217, 8'd204, 8'd102};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd212, 8'd171, 8'd43};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd240, 8'd168, 8'd34};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd238, 8'd152, 8'd33};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd230, 8'd136, 8'd23};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd219, 8'd113, 8'd11};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd214, 8'd99, 8'd6};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd217, 8'd97, 8'd10};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd223, 8'd105, 8'd17};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd228, 8'd113, 8'd22};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd230, 8'd117, 8'd23};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd210, 8'd108, 8'd10};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd206, 8'd95, 8'd6};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd214, 8'd96, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd168, 8'd61, 8'd7};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd142, 8'd56, 8'd5};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd232, 8'd169, 8'd98};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd251, 8'd199, 8'd97};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd196, 8'd147, 8'd19};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd235, 8'd173, 8'd88};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd241, 8'd193, 8'd93};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd239, 8'd191, 8'd83};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd201, 8'd122, 8'd29};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd205, 8'd94, 8'd25};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd149, 8'd45, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd211, 8'd161, 8'd76};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd221, 8'd223, 8'd114};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd243, 8'd212, 8'd129};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd168, 8'd78, 8'd26};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd146, 8'd73, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd179};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd170};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd152};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd228, 8'd160, 8'd79};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd235, 8'd130, 8'd47};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd239, 8'd138, 8'd70};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd215, 8'd121, 8'd51};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd218, 8'd126, 8'd53};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd229, 8'd134, 8'd52};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd226, 8'd124, 8'd42};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd208, 8'd107, 8'd39};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd153, 8'd66, 8'd21};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd166, 8'd94, 8'd69};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd246, 8'd212, 8'd141};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd175};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd231, 8'd189, 8'd139};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd214, 8'd161, 8'd91};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd212, 8'd146, 8'd86};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd163, 8'd94, 8'd65};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd240, 8'd190, 8'd165};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd188};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd133};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd185, 8'd132, 8'd38};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd222, 8'd145, 8'd55};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd206, 8'd116, 8'd38};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd159, 8'd76, 8'd8};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd189, 8'd121, 8'd50};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd111};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd108};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd241, 8'd162, 8'd96};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd140, 8'd55, 8'd0};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd189, 8'd130, 8'd52};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd254, 8'd235, 8'd140};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd228, 8'd209, 8'd114};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd172, 8'd110, 8'd33};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd152, 8'd64, 8'd0};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd218, 8'd137, 8'd72};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd108};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd251, 8'd205, 8'd107};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd226, 8'd178, 8'd78};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd219, 8'd152, 8'd63};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd238, 8'd146, 8'd79};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd212, 8'd124, 8'd78};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd160, 8'd101, 8'd67};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd208};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd191};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd169};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd215, 8'd157, 8'd94};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd240, 8'd162, 8'd90};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd225, 8'd132, 8'd52};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd237, 8'd142, 8'd52};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd225, 8'd131, 8'd35};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd217, 8'd128, 8'd28};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd216, 8'd116, 8'd20};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd215, 8'd121, 8'd21};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd228, 8'd141, 8'd28};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd231, 8'd144, 8'd15};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd240, 8'd158, 8'd20};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd228, 8'd161, 8'd28};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd204, 8'd164, 8'd50};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd238, 8'd220, 8'd120};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd212, 8'd169};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd236, 8'd128, 8'd27};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd252, 8'd155, 8'd24};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd241, 8'd156, 8'd50};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd214, 8'd98, 8'd49};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd206, 8'd47, 8'd43};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd209, 8'd29, 8'd38};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd206, 8'd34, 8'd32};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd207, 8'd33, 8'd32};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd207, 8'd31, 8'd31};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd207, 8'd28, 8'd31};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd203, 8'd27, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd197, 8'd24, 8'd26};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd192, 8'd23, 8'd26};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd187, 8'd23, 8'd24};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd146, 8'd10, 8'd24};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd228, 8'd118, 8'd121};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd185};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd136: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd187, 8'd133, 8'd121};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd145, 8'd45, 8'd45};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd145, 8'd0, 8'd2};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd184, 8'd0, 8'd13};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd199, 8'd20, 8'd26};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd193, 8'd28, 8'd24};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd193, 8'd28, 8'd22};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd195, 8'd23, 8'd19};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd209, 8'd30, 8'd36};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd200, 8'd29, 8'd21};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd199, 8'd29, 8'd14};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd226, 8'd36, 8'd38};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd223, 8'd14, 8'd36};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd224, 8'd25, 8'd32};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd209, 8'd54, 8'd10};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd252, 8'd137, 8'd46};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd242, 8'd145, 8'd42};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd235, 8'd140, 8'd22};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd245, 8'd176, 8'd119};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd238, 8'd215, 8'd161};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd217, 8'd182, 8'd88};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd207, 8'd165, 8'd47};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd179, 8'd41};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd239, 8'd157, 8'd19};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd229, 8'd136, 8'd7};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd231, 8'd125, 8'd16};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd227, 8'd113, 8'd25};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd216, 8'd104, 8'd20};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd211, 8'd107, 8'd10};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd215, 8'd118, 8'd5};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd216, 8'd101, 8'd12};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd226, 8'd106, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd217, 8'd97, 8'd37};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd188, 8'd73, 8'd19};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd142, 8'd43, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd217, 8'd142, 8'd51};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd236, 8'd186, 8'd63};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd233, 8'd198, 8'd54};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd237, 8'd198, 8'd107};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd247, 8'd196, 8'd91};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd220, 8'd146, 8'd41};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd225, 8'd129, 8'd53};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd193, 8'd87, 8'd47};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd119, 8'd23, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd234, 8'd162, 8'd80};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd252, 8'd201, 8'd74};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd130};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd169, 8'd95, 8'd20};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd152, 8'd57, 8'd0};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd84};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd255, 8'd226, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd246, 8'd224, 8'd113};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd236, 8'd196, 8'd75};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd221, 8'd155, 8'd33};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd175, 8'd110, 8'd10};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd177, 8'd105, 8'd7};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd230, 8'd149, 8'd57};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd218, 8'd126, 8'd41};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd210, 8'd108, 8'd33};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd217, 8'd109, 8'd45};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd179, 8'd68, 8'd13};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd199, 8'd87, 8'd37};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd250, 8'd204, 8'd108};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd105};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd229, 8'd162, 8'd71};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd218, 8'd140, 8'd57};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd219, 8'd138, 8'd59};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd189, 8'd111, 8'd39};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd204, 8'd133, 8'd67};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd156};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd208, 8'd80};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd235, 8'd175, 8'd51};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd184, 8'd123, 8'd6};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd155, 8'd93, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd182, 8'd118, 8'd18};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd237, 8'd172, 8'd80};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd114};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd255, 8'd194, 8'd113};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd214, 8'd122, 8'd81};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd162, 8'd83, 8'd14};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd201, 8'd139, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd251, 8'd199, 8'd63};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd237, 8'd185, 8'd49};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd198, 8'd136, 8'd27};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd172, 8'd93, 8'd24};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd182, 8'd90, 8'd49};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd190, 8'd105};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd250, 8'd191, 8'd97};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd240, 8'd190, 8'd91};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd219, 8'd148, 8'd60};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd255, 8'd158, 8'd92};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd223, 8'd118, 8'd73};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd145, 8'd80, 8'd40};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd232, 8'd191};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd207};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd180};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd224, 8'd158, 8'd100};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd244, 8'd160, 8'd87};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd222, 8'd136, 8'd49};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd210, 8'd123, 8'd28};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd222, 8'd131, 8'd38};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd228, 8'd128, 8'd40};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd196, 8'd120, 8'd10};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd222, 8'd148, 8'd15};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd229, 8'd160, 8'd20};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd230, 8'd166, 8'd34};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd221, 8'd175, 8'd27};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd197, 8'd173, 8'd15};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd213, 8'd198, 8'd95};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd177};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd225, 8'd131, 8'd18};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd234, 8'd145, 8'd17};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd247, 8'd160, 8'd47};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd227, 8'd102, 8'd22};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd199, 8'd25, 8'd26};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd225, 8'd39, 8'd40};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd218, 8'd30, 8'd29};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd210, 8'd25, 8'd23};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd205, 8'd23, 8'd19};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd213, 8'd38, 8'd33};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd194, 8'd24, 8'd24};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd177, 8'd13, 8'd22};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd188, 8'd29, 8'd47};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd173, 8'd17, 8'd39};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd199, 8'd164, 8'd170};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd250, 8'd224, 8'd227};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd137: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd218, 8'd139, 8'd134};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd162, 8'd44, 8'd44};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd175, 8'd22, 8'd25};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd192, 8'd19, 8'd23};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd195, 8'd16, 8'd19};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd210, 8'd34, 8'd34};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd202, 8'd27, 8'd34};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd206, 8'd42, 8'd32};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd204, 8'd43, 8'd25};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd211, 8'd37, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd205, 8'd17, 8'd32};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd209, 8'd29, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd203, 8'd61, 8'd13};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd252, 8'd145, 8'd51};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd243, 8'd146, 8'd41};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd235, 8'd140, 8'd20};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd244, 8'd175, 8'd116};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd255, 8'd245, 8'd202};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd239, 8'd211, 8'd137};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd212, 8'd178, 8'd81};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd232, 8'd165, 8'd35};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd237, 8'd163, 8'd28};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd239, 8'd153, 8'd18};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd233, 8'd135, 8'd12};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd224, 8'd117, 8'd13};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd217, 8'd110, 8'd16};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd213, 8'd109, 8'd10};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd209, 8'd111, 8'd4};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd213, 8'd102, 8'd10};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd244, 8'd129, 8'd48};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd210, 8'd90, 8'd27};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd198, 8'd83, 8'd28};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd156, 8'd54, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd164, 8'd82, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd254, 8'd194, 8'd80};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd245, 8'd198, 8'd66};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd240, 8'd195, 8'd104};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd246, 8'd189, 8'd84};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd223, 8'd146, 8'd42};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd220, 8'd123, 8'd46};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd196, 8'd89, 8'd45};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd139, 8'd42, 8'd0};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd237, 8'd163, 8'd78};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd73};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd255, 8'd207, 8'd113};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd186, 8'd108, 8'd26};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd171, 8'd72, 8'd4};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd180, 8'd96, 8'd23};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd194, 8'd144, 8'd55};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd230, 8'd197, 8'd90};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd255, 8'd206, 8'd93};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd255, 8'd200, 8'd85};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd255, 8'd201, 8'd102};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd248, 8'd185, 8'd88};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd255, 8'd195, 8'd100};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd234, 8'd153, 8'd62};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd209, 8'd118, 8'd37};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd203, 8'd107, 8'd33};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd173, 8'd75, 8'd10};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd188, 8'd90, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd251, 8'd197, 8'd99};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd196, 8'd101};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd236, 8'd163, 8'd69};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd216, 8'd135, 8'd44};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd212, 8'd128, 8'd42};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd186, 8'd105, 8'd24};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd180, 8'd107, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd217, 8'd149, 8'd74};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd251, 8'd197, 8'd75};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd255, 8'd202, 8'd83};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd252, 8'd197, 8'd81};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd244, 8'd188, 8'd79};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd253, 8'd195, 8'd95};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd255, 8'd205, 8'd111};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd250, 8'd191, 8'd101};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd222, 8'd162, 8'd74};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd214, 8'd122, 8'd71};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd170, 8'd88, 8'd14};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd205, 8'd136, 8'd32};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd252, 8'd194, 8'd68};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd245, 8'd187, 8'd61};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd214, 8'd145, 8'd41};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd182, 8'd100, 8'd26};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd176, 8'd84, 8'd33};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd243, 8'd176, 8'd89};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd246, 8'd196, 8'd101};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd250, 8'd207, 8'd105};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd220, 8'd155, 8'd63};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd227, 8'd133, 8'd59};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd187, 8'd91, 8'd33};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd142, 8'd81, 8'd26};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd229, 8'd172};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd255, 8'd235, 8'd180};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd247, 8'd202, 8'd145};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd204, 8'd130, 8'd65};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd226, 8'd139, 8'd60};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd222, 8'd133, 8'd41};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd216, 8'd130, 8'd31};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd221, 8'd131, 8'd34};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd215, 8'd118, 8'd24};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd217, 8'd138, 8'd35};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd218, 8'd142, 8'd32};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd235, 8'd167, 8'd32};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd230, 8'd176, 8'd15};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd204, 8'd165, 8'd10};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd218, 8'd191, 8'd84};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd252, 8'd234, 8'd188};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd174};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd225, 8'd131, 8'd17};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd235, 8'd146, 8'd18};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd250, 8'd163, 8'd50};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd232, 8'd107, 8'd27};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd199, 8'd27, 8'd27};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd221, 8'd37, 8'd37};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd206, 8'd46, 8'd34};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd194, 8'd23, 8'd15};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd209, 8'd25, 8'd23};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd192, 8'd6, 8'd9};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd184, 8'd11, 8'd17};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd161, 8'd17, 8'd26};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd153, 8'd44, 8'd50};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd248, 8'd161, 8'd169};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd245, 8'd216, 8'd220};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd138: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd227, 8'd187, 8'd175};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd175, 8'd69, 8'd69};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd170, 8'd6, 8'd15};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd193, 8'd9, 8'd19};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd189, 8'd6, 8'd11};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd186, 8'd15, 8'd23};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd194, 8'd33, 8'd25};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd195, 8'd40, 8'd22};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd201, 8'd42, 8'd36};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd205, 8'd38, 8'd46};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd202, 8'd45, 8'd38};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd199, 8'd69, 8'd17};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd152, 8'd57};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd245, 8'd149, 8'd39};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd235, 8'd141, 8'd17};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd241, 8'd173, 8'd112};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd192};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd234, 8'd213, 8'd150};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd220, 8'd166, 8'd57};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd226, 8'd165, 8'd40};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd234, 8'd163, 8'd21};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd237, 8'd152, 8'd10};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd229, 8'd134, 8'd8};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd217, 8'd116, 8'd8};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd209, 8'd110, 8'd8};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd207, 8'd110, 8'd7};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd100, 8'd2};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd230, 8'd120, 8'd33};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd206, 8'd92, 8'd21};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd206, 8'd92, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd186, 8'd81, 8'd16};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd154, 8'd61, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd255, 8'd183, 8'd83};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd254, 8'd187, 8'd74};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd233, 8'd178, 8'd85};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd240, 8'd175, 8'd73};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd231, 8'd149, 8'd47};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd222, 8'd125, 8'd46};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd210, 8'd105, 8'd50};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd174, 8'd78, 8'd20};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd238, 8'd158, 8'd69};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd246, 8'd182, 8'd59};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd248, 8'd185, 8'd80};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd211, 8'd126, 8'd35};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd220, 8'd119, 8'd39};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd183, 8'd94, 8'd12};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd165, 8'd101, 8'd11};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd207, 8'd158, 8'd55};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd232, 8'd169, 8'd63};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd255, 8'd182, 8'd76};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd255, 8'd203, 8'd107};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd255, 8'd198, 8'd101};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd255, 8'd199, 8'd103};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd245, 8'd171, 8'd76};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd220, 8'd139, 8'd48};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd202, 8'd118, 8'd32};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd179, 8'd94, 8'd13};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd181, 8'd95, 8'd18};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd250, 8'd184, 8'd87};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd191, 8'd93};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd251, 8'd171, 8'd72};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd234, 8'd148, 8'd49};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd229, 8'd141, 8'd43};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd214, 8'd130, 8'd32};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd192, 8'd113, 8'd18};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd182, 8'd109, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd205, 8'd154, 8'd39};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd230, 8'd178, 8'd66};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd250, 8'd198, 8'd88};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd252, 8'd199, 8'd93};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd251, 8'd197, 8'd97};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd248, 8'd194, 8'd98};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd230, 8'd175, 8'd82};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd207, 8'd152, 8'd61};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd219, 8'd126, 8'd57};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd188, 8'd103, 8'd22};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd215, 8'd139, 8'd43};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd253, 8'd185, 8'd76};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd252, 8'd184, 8'd75};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd231, 8'd155, 8'd59};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd199, 8'd114, 8'd33};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd181, 8'd88, 8'd19};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd228, 8'd168, 8'd82};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd237, 8'd191, 8'd97};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd245, 8'd206, 8'd105};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd234, 8'd176, 8'd79};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd238, 8'd154, 8'd68};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd206, 8'd119, 8'd42};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd172, 8'd110, 8'd35};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd232, 8'd199, 8'd120};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd246, 8'd207, 8'd138};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd243, 8'd183, 8'd111};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd214, 8'd131, 8'd53};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd235, 8'd141, 8'd53};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd233, 8'd144, 8'd44};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd226, 8'd141, 8'd35};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd226, 8'd139, 8'd34};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd215, 8'd121, 8'd21};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd50};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd229, 8'd154, 8'd52};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd230, 8'd171, 8'd33};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd216, 8'd176, 8'd0};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd208, 8'd181, 8'd42};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd245, 8'd221, 8'd175};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd254, 8'd194, 8'd168};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd225, 8'd130, 8'd14};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd237, 8'd148, 8'd18};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd253, 8'd166, 8'd53};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd238, 8'd115, 8'd35};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd199, 8'd29, 8'd29};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd215, 8'd33, 8'd32};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd185, 8'd44, 8'd24};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd204, 8'd44, 8'd32};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd192, 8'd8, 8'd8};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd202, 8'd15, 8'd24};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd173, 8'd11, 8'd24};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd149, 8'd40, 8'd46};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd215, 8'd167, 8'd163};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd139: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd238, 8'd187, 8'd183};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd189, 8'd74, 8'd79};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd173, 8'd9, 8'd20};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd205, 8'd19, 8'd32};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd190, 8'd18, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd186, 8'd21, 8'd17};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd186, 8'd24, 8'd13};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd196, 8'd34, 8'd31};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd208, 8'd49, 8'd54};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd194, 8'd46, 8'd36};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd194, 8'd67, 8'd12};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd56};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd248, 8'd152, 8'd39};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd234, 8'd141, 8'd12};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd238, 8'd170, 8'd105};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd235, 8'd197, 8'd116};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd213, 8'd169, 8'd60};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd212, 8'd156, 8'd17};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd233, 8'd164, 8'd11};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd240, 8'd157, 8'd15};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd222, 8'd130, 8'd7};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd208, 8'd113, 8'd5};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd212, 8'd116, 8'd13};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd215, 8'd116, 8'd12};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd202, 8'd99, 8'd4};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd216, 8'd109, 8'd27};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd202, 8'd91, 8'd19};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd198, 8'd89, 8'd20};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd174, 8'd73, 8'd0};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd203, 8'd112, 8'd23};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd202, 8'd115, 8'd18};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd207, 8'd141, 8'd45};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd218, 8'd145, 8'd43};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd228, 8'd142, 8'd43};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd220, 8'd124, 8'd38};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd218, 8'd117, 8'd47};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd197, 8'd103, 8'd29};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd221, 8'd139, 8'd40};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd216, 8'd144, 8'd23};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd224, 8'd149, 8'd34};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd213, 8'd124, 8'd20};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd242, 8'd142, 8'd48};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd223, 8'd130, 8'd37};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd189, 8'd113, 8'd17};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd189, 8'd121, 8'd20};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd189, 8'd111, 8'd11};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd209, 8'd120, 8'd20};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd188, 8'd124, 8'd34};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd203, 8'd137, 8'd43};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd219, 8'd146, 8'd51};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd227, 8'd149, 8'd51};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd220, 8'd137, 8'd41};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd205, 8'd121, 8'd25};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd195, 8'd112, 8'd20};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd188, 8'd104, 8'd14};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd204, 8'd129, 8'd28};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd221, 8'd142, 8'd41};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd231, 8'd148, 8'd42};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd233, 8'd147, 8'd36};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd239, 8'd152, 8'd39};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd244, 8'd160, 8'd48};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd230, 8'd150, 8'd39};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd206, 8'd130, 8'd18};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd187, 8'd129, 8'd22};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd200, 8'd142, 8'd35};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd206, 8'd147, 8'd43};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd202, 8'd143, 8'd41};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd205, 8'd145, 8'd47};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd217, 8'd157, 8'd61};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd227, 8'd166, 8'd73};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd227, 8'd166, 8'd73};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd241, 8'd151, 8'd65};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd211, 8'd126, 8'd36};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd207, 8'd126, 8'd34};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd213, 8'd137, 8'd41};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd212, 8'd136, 8'd40};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd217, 8'd136, 8'd44};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd220, 8'd135, 8'd45};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd216, 8'd126, 8'd40};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd201, 8'd140, 8'd59};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd201, 8'd150, 8'd61};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd206, 8'd157, 8'd62};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd217, 8'd154, 8'd57};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd233, 8'd154, 8'd62};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd222, 8'd138, 8'd50};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd193, 8'd123, 8'd35};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd199, 8'd145, 8'd55};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd196, 8'd141, 8'd58};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd216, 8'd144, 8'd60};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd220, 8'd128, 8'd41};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd236, 8'd139, 8'd44};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd226, 8'd139, 8'd33};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd217, 8'd137, 8'd24};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd229, 8'd147, 8'd35};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd231, 8'd145, 8'd36};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd234, 8'd160, 8'd37};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd241, 8'd176, 8'd46};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd217, 8'd170, 8'd22};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd206, 8'd175, 8'd33};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd239, 8'd218, 8'd135};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd249, 8'd188, 8'd159};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd227, 8'd130, 8'd13};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd239, 8'd151, 8'd18};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd53};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd242, 8'd121, 8'd40};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd197, 8'd29, 8'd29};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd207, 8'd27, 8'd28};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd198, 8'd40, 8'd28};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd196, 8'd29, 8'd23};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd205, 8'd32, 8'd34};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd172, 8'd10, 8'd21};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd169, 8'd43, 8'd54};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd233, 8'd164, 8'd167};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd140: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd239, 8'd188, 8'd184};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd196, 8'd81, 8'd88};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd167, 8'd5, 8'd20};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd188, 8'd23, 8'd37};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd192, 8'd22, 8'd23};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd202, 8'd24, 8'd20};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd197, 8'd18, 8'd22};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd199, 8'd29, 8'd40};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd184, 8'd33, 8'd24};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd201, 8'd67, 8'd14};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd146, 8'd55};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd251, 8'd156, 8'd36};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd234, 8'd142, 8'd9};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd235, 8'd168, 8'd98};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd184};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd219, 8'd191, 8'd108};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd199, 8'd159, 8'd35};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd218, 8'd162, 8'd13};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd239, 8'd167, 8'd21};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd236, 8'd152, 8'd20};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd220, 8'd131, 8'd13};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd213, 8'd121, 8'd10};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd214, 8'd122, 8'd13};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd197, 8'd101, 8'd0};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd223, 8'd123, 8'd29};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd210, 8'd106, 8'd19};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd209, 8'd104, 8'd21};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd213, 8'd111, 8'd27};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd191, 8'd91, 8'd3};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd189, 8'd91, 8'd0};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd209, 8'd134, 8'd33};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd219, 8'd140, 8'd39};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd232, 8'd146, 8'd47};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd223, 8'd132, 8'd39};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd228, 8'd136, 8'd49};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd222, 8'd133, 8'd41};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd220, 8'd137, 8'd31};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd214, 8'd138, 8'd18};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd227, 8'd144, 8'd22};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd225, 8'd138, 8'd22};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd236, 8'd144, 8'd35};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd242, 8'd151, 8'd46};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd224, 8'd141, 8'd37};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd208, 8'd129, 8'd26};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd209, 8'd126, 8'd24};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd211, 8'd122, 8'd22};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd199, 8'd119, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd212, 8'd129, 8'd37};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd216, 8'd129, 8'd34};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd226, 8'd136, 8'd39};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd228, 8'd136, 8'd37};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd222, 8'd130, 8'd31};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd225, 8'd137, 8'd39};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd220, 8'd133, 8'd36};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd204, 8'd122, 8'd20};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd213, 8'd132, 8'd25};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd231, 8'd147, 8'd35};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd238, 8'd155, 8'd37};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd237, 8'd154, 8'd34};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd240, 8'd160, 8'd37};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd236, 8'd160, 8'd38};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd222, 8'd148, 8'd27};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd218, 8'd147, 8'd43};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd218, 8'd146, 8'd44};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd214, 8'd142, 8'd42};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd210, 8'd138, 8'd40};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd216, 8'd143, 8'd48};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd229, 8'd156, 8'd62};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd239, 8'd166, 8'd74};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd242, 8'd168, 8'd79};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd245, 8'd162, 8'd66};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd234, 8'd154, 8'd59};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd226, 8'd147, 8'd54};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd220, 8'd143, 8'd51};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd214, 8'd137, 8'd45};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd223, 8'd144, 8'd51};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd238, 8'd158, 8'd63};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd240, 8'd157, 8'd61};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd228, 8'd161, 8'd80};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd224, 8'd162, 8'd77};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd230, 8'd169, 8'd80};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd237, 8'd170, 8'd79};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd243, 8'd166, 8'd76};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd247, 8'd166, 8'd77};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd242, 8'd165, 8'd77};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd235, 8'd164, 8'd74};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd202, 8'd138, 8'd48};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd224, 8'd147, 8'd55};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd234, 8'd143, 8'd50};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd229, 8'd137, 8'd36};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd214, 8'd134, 8'd23};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd205, 8'd133, 8'd15};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd228, 8'd153, 8'd34};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd240, 8'd159, 8'd42};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd235, 8'd174, 8'd24};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd226, 8'd179, 8'd11};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd208, 8'd176, 8'd29};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd224, 8'd201, 8'd125};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd228};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd243, 8'd180, 8'd147};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd229, 8'd133, 8'd13};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd241, 8'd153, 8'd19};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd253, 8'd168, 8'd52};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd244, 8'd123, 8'd42};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd192, 8'd26, 8'd26};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd200, 8'd22, 8'd22};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd205, 8'd17, 8'd18};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd200, 8'd26, 8'd28};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd168, 8'd22, 8'd25};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd147, 8'd37, 8'd40};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd213, 8'd142, 8'd146};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd141: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd240, 8'd180, 8'd179};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd164, 8'd57, 8'd63};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd152, 8'd15, 8'd22};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd176, 8'd16, 8'd18};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd219, 8'd31, 8'd32};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd212, 8'd16, 8'd28};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd201, 8'd20, 8'd35};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd188, 8'd34, 8'd26};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd216, 8'd85, 8'd31};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd151, 8'd57};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd254, 8'd160, 8'd36};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd234, 8'd143, 8'd3};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd232, 8'd166, 8'd92};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd255, 8'd252, 8'd234};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd239, 8'd226, 8'd173};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd215, 8'd187, 8'd88};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd206, 8'd162, 8'd31};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd225, 8'd161, 8'd25};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd247, 8'd170, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd238, 8'd155, 8'd27};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd215, 8'd130, 8'd3};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd197, 8'd107, 8'd0};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd207, 8'd117, 8'd7};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd207, 8'd114, 8'd10};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd215, 8'd119, 8'd17};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd210, 8'd112, 8'd13};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd223, 8'd125, 8'd28};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd220, 8'd121, 8'd27};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd215, 8'd116, 8'd22};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd225, 8'd144, 8'd37};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd230, 8'd148, 8'd46};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd229, 8'd145, 8'd46};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd221, 8'd137, 8'd38};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd228, 8'd145, 8'd41};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd230, 8'd148, 8'd38};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd224, 8'd145, 8'd27};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd227, 8'd148, 8'd29};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd238, 8'd156, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd243, 8'd161, 8'd35};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd230, 8'd147, 8'd25};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd228, 8'd145, 8'd27};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd229, 8'd145, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd233, 8'd148, 8'd39};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd241, 8'd156, 8'd49};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd226, 8'd141, 8'd35};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd227, 8'd140, 8'd47};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd231, 8'd141, 8'd45};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd230, 8'd138, 8'd39};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd234, 8'd138, 8'd36};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd234, 8'd138, 8'd35};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd229, 8'd137, 8'd34};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd231, 8'd144, 8'd41};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd229, 8'd143, 8'd44};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd225, 8'd146, 8'd41};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd229, 8'd151, 8'd42};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd238, 8'd161, 8'd45};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd240, 8'd164, 8'd44};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd231, 8'd157, 8'd32};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd226, 8'd155, 8'd29};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd227, 8'd157, 8'd33};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd226, 8'd156, 8'd34};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd230, 8'd160, 8'd48};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd228, 8'd158, 8'd47};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd228, 8'd157, 8'd49};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd233, 8'd162, 8'd58};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd71};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd245, 8'd172, 8'd78};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd243, 8'd170, 8'd78};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd239, 8'd165, 8'd76};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd234, 8'd162, 8'd62};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd243, 8'd171, 8'd71};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd240, 8'd168, 8'd68};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd237, 8'd168, 8'd67};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd230, 8'd161, 8'd60};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd230, 8'd158, 8'd58};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd243, 8'd171, 8'd71};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd242, 8'd170, 8'd70};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd235, 8'd169, 8'd85};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd230, 8'd165, 8'd81};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd242, 8'd178, 8'd91};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd241, 8'd179, 8'd94};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd235, 8'd173, 8'd88};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd244, 8'd178, 8'd94};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd244, 8'd173, 8'd91};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd238, 8'd162, 8'd84};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd235, 8'd174, 8'd81};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd240, 8'd167, 8'd75};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd240, 8'd155, 8'd62};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd218, 8'd134, 8'd35};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd214, 8'd142, 8'd31};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd214, 8'd152, 8'd31};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd239, 8'd173, 8'd50};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd247, 8'd176, 8'd52};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd235, 8'd187, 8'd29};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd205, 8'd170, 8'd8};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd220, 8'd198, 8'd86};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd255, 8'd240, 8'd219};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd236, 8'd172, 8'd137};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd234, 8'd135, 8'd15};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd246, 8'd155, 8'd22};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd248, 8'd163, 8'd47};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd239, 8'd120, 8'd38};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd186, 8'd22, 8'd23};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd194, 8'd18, 8'd20};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd190, 8'd3, 8'd14};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd173, 8'd16, 8'd23};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd143, 8'd34, 8'd37};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd207, 8'd147, 8'd146};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd142: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd246, 8'd226, 8'd219};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd206};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd166, 8'd66, 8'd64};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd157, 8'd19, 8'd16};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd205, 8'd21, 8'd23};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd218, 8'd16, 8'd32};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd210, 8'd25, 8'd43};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd185, 8'd34, 8'd25};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd215, 8'd96, 8'd38};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd161, 8'd62};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd255, 8'd163, 8'd34};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd234, 8'd143, 8'd2};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd229, 8'd163, 8'd85};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd244, 8'd226, 8'd154};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd217, 8'd179, 8'd72};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd216, 8'd158, 8'd35};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd239, 8'd166, 8'd38};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd246, 8'd165, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd233, 8'd150, 8'd8};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd207, 8'd117, 8'd7};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd218, 8'd131, 8'd18};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd200, 8'd113, 8'd0};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd206, 8'd119, 8'd4};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd201, 8'd111, 8'd0};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd203, 8'd113, 8'd1};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd213, 8'd120, 8'd14};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd212, 8'd116, 8'd13};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd226, 8'd141, 8'd32};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd229, 8'd148, 8'd43};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd216, 8'd137, 8'd36};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd215, 8'd138, 8'd32};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd220, 8'd148, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd220, 8'd146, 8'd21};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd214, 8'd139, 8'd14};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd225, 8'd146, 8'd27};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd227, 8'd148, 8'd19};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd230, 8'd157, 8'd26};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd227, 8'd159, 8'd26};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd212, 8'd139, 8'd10};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd219, 8'd136, 8'd14};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd235, 8'd150, 8'd33};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd227, 8'd146, 8'd29};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd217, 8'd142, 8'd27};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd213, 8'd131, 8'd29};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd213, 8'd130, 8'd24};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd222, 8'd135, 8'd29};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd223, 8'd137, 8'd26};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd225, 8'd139, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd223, 8'd141, 8'd33};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd213, 8'd136, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd210, 8'd135, 8'd33};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd214, 8'd137, 8'd29};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd222, 8'd149, 8'd36};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd224, 8'd155, 8'd36};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd222, 8'd156, 8'd33};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd226, 8'd162, 8'd38};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd229, 8'd167, 8'd44};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd232, 8'd170, 8'd49};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd235, 8'd172, 8'd56};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd224, 8'd166, 8'd40};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd222, 8'd164, 8'd39};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd225, 8'd166, 8'd46};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd233, 8'd173, 8'd59};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd239, 8'd178, 8'd72};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd238, 8'd176, 8'd77};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd236, 8'd173, 8'd78};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd235, 8'd171, 8'd81};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd235, 8'd175, 8'd77};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd76};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd216, 8'd155, 8'd48};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd212, 8'd150, 8'd39};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd211, 8'd149, 8'd38};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd214, 8'd153, 8'd46};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd239, 8'd177, 8'd76};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd243, 8'd183, 8'd85};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd234, 8'd181, 8'd87};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd221, 8'd167, 8'd77};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd239, 8'd187, 8'd101};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd235, 8'd190, 8'd105};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd228, 8'd191, 8'd110};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd241, 8'd202, 8'd123};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd237, 8'd187, 8'd114};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd238, 8'd178, 8'd108};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd223, 8'd169, 8'd79};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd221, 8'd155, 8'd68};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd225, 8'd149, 8'd61};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd204, 8'd132, 8'd34};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd218, 8'd158, 8'd48};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd229, 8'd175, 8'd53};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd251, 8'd194, 8'd65};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd251, 8'd186, 8'd56};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd223, 8'd182, 8'd40};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd218, 8'd187, 8'd79};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd243, 8'd226, 8'd174};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd230, 8'd165, 8'd127};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd238, 8'd140, 8'd17};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd247, 8'd157, 8'd21};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd242, 8'd157, 8'd40};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd233, 8'd114, 8'd32};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd180, 8'd16, 8'd17};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd190, 8'd16, 8'd17};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd173, 8'd28, 8'd35};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd149, 8'd33, 8'd36};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd221, 8'd151, 8'd151};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd143: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd229, 8'd251, 8'd228};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd238, 8'd170, 8'd159};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd161, 8'd44, 8'd34};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd177, 8'd1, 8'd3};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd207, 8'd5, 8'd21};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd201, 8'd18, 8'd36};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd160, 8'd18, 8'd6};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd196, 8'd88, 8'd24};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd168, 8'd64};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd255, 8'd164, 8'd33};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd234, 8'd143, 8'd0};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd228, 8'd163, 8'd83};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd255, 8'd250, 8'd195};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd238, 8'd201, 8'd112};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd215, 8'd159, 8'd48};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd222, 8'd151, 8'd27};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd240, 8'd163, 8'd21};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd252, 8'd173, 8'd20};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd236, 8'd146, 8'd36};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd224, 8'd137, 8'd24};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd220, 8'd135, 8'd16};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd217, 8'd135, 8'd10};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd224, 8'd142, 8'd17};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd231, 8'd146, 8'd27};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd226, 8'd136, 8'd22};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd236, 8'd144, 8'd33};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd240, 8'd156, 8'd42};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd249, 8'd168, 8'd61};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd233, 8'd155, 8'd54};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd241, 8'd169, 8'd59};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd244, 8'd176, 8'd51};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd235, 8'd167, 8'd34};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd228, 8'd155, 8'd27};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd237, 8'd161, 8'd41};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd230, 8'd153, 8'd23};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd225, 8'd157, 8'd24};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd247, 8'd185, 8'd48};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd230, 8'd164, 8'd28};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd237, 8'd158, 8'd31};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd255, 8'd172, 8'd48};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd232, 8'd153, 8'd32};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd242, 8'd172, 8'd50};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd227, 8'd155, 8'd44};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd222, 8'd149, 8'd36};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd234, 8'd159, 8'd44};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd233, 8'd156, 8'd40};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd236, 8'd161, 8'd46};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd239, 8'd169, 8'd57};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd223, 8'd159, 8'd51};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd225, 8'd162, 8'd56};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd239, 8'd167, 8'd57};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd251, 8'd181, 8'd67};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd243, 8'd178, 8'd60};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd230, 8'd170, 8'd48};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd235, 8'd179, 8'd56};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd242, 8'd186, 8'd65};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd236, 8'd179, 8'd63};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd234, 8'd174, 8'd62};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd232, 8'd189, 8'd50};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd230, 8'd186, 8'd51};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd232, 8'd188, 8'd57};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd236, 8'd190, 8'd68};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd233, 8'd185, 8'd74};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd228, 8'd179, 8'd74};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd227, 8'd177, 8'd78};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd231, 8'd181, 8'd86};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd233, 8'd180, 8'd84};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd241, 8'd188, 8'd84};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd228, 8'd175, 8'd61};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd239, 8'd185, 8'd63};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd246, 8'd192, 8'd70};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd237, 8'd184, 8'd70};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd243, 8'd190, 8'd86};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd236, 8'd183, 8'd87};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd240, 8'd201, 8'd100};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd224, 8'd184, 8'd88};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd245, 8'd205, 8'd117};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd229, 8'd201, 8'd117};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd217, 8'd202, 8'd121};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd239, 8'd223, 8'd146};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd249, 8'd218, 8'd151};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd167};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd240, 8'd192, 8'd107};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd244, 8'd183, 8'd100};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd254, 8'd184, 8'd98};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd226, 8'd160, 8'd64};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd232, 8'd178, 8'd69};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd231, 8'd182, 8'd61};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd238, 8'd185, 8'd55};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd231, 8'd168, 8'd37};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd204, 8'd168, 8'd46};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd252, 8'd219, 8'd166};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd226, 8'd161, 8'd123};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd241, 8'd141, 8'd17};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd248, 8'd158, 8'd22};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd238, 8'd153, 8'd36};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd227, 8'd111, 8'd28};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd176, 8'd13, 8'd14};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd189, 8'd15, 8'd16};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd139, 8'd39, 8'd37};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd233, 8'd154, 8'd150};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd144: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd213, 8'd174, 8'd157};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd161, 8'd71, 8'd63};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd155, 8'd1, 8'd13};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd209, 8'd12, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd210, 8'd23, 8'd16};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd181, 8'd51, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd249, 8'd170, 8'd67};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd252, 8'd147, 8'd38};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd245, 8'd153, 8'd44};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd213, 8'd144, 8'd67};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd199};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd221, 8'd213, 8'd150};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd195, 8'd162, 8'd57};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd208, 8'd147, 8'd5};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd242, 8'd163, 8'd0};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd221, 8'd162, 8'd6};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd220, 8'd164, 8'd9};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd221, 8'd166, 8'd14};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd222, 8'd168, 8'd20};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd223, 8'd170, 8'd28};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd225, 8'd173, 8'd37};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd224, 8'd174, 8'd41};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd224, 8'd175, 8'd44};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd231, 8'd168, 8'd62};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd248, 8'd185, 8'd79};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd243, 8'd181, 8'd72};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd238, 8'd176, 8'd65};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd248, 8'd186, 8'd73};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd242, 8'd181, 8'd66};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd236, 8'd175, 8'd58};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd252, 8'd192, 8'd72};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd245, 8'd185, 8'd65};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd247, 8'd188, 8'd68};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd245, 8'd193, 8'd73};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd246, 8'd195, 8'd77};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd245, 8'd196, 8'd78};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd246, 8'd195, 8'd80};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd248, 8'd195, 8'd83};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd251, 8'd195, 8'd84};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd240, 8'd194, 8'd82};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd239, 8'd193, 8'd81};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd240, 8'd194, 8'd82};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd244, 8'd198, 8'd86};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd248, 8'd202, 8'd90};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd252, 8'd204, 8'd93};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd251, 8'd203, 8'd92};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd249, 8'd201, 8'd90};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd246, 8'd204, 8'd86};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd255, 8'd214, 8'd96};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd250, 8'd209, 8'd93};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd249, 8'd208, 8'd94};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd106};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd106};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd252, 8'd215, 8'd101};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd113};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd255, 8'd233, 8'd123};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd250, 8'd219, 8'd111};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd253, 8'd220, 8'd115};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd255, 8'd225, 8'd125};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd255, 8'd222, 8'd127};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd139};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd145};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd245, 8'd224, 8'd133};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd253, 8'd223, 8'd151};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd253, 8'd221, 8'd146};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd255, 8'd227, 8'd146};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd253, 8'd221, 8'd138};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd235, 8'd203, 8'd120};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd247, 8'd214, 8'd137};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd255, 8'd238, 8'd167};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd255, 8'd243, 8'd178};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd255, 8'd230, 8'd168};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd255, 8'd231, 8'd173};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd255, 8'd234, 8'd181};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd255, 8'd236, 8'd190};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd255, 8'd239, 8'd200};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd255, 8'd242, 8'd209};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd255, 8'd244, 8'd216};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd255, 8'd246, 8'd221};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd250, 8'd229, 8'd182};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd248, 8'd220, 8'd155};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd248, 8'd212, 8'd118};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd250, 8'd208, 8'd88};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd252, 8'd206, 8'd71};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd241, 8'd198, 8'd60};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd222, 8'd183, 8'd54};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd207, 8'd171, 8'd49};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd250, 8'd234, 8'd174};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd252, 8'd239, 8'd197};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd255, 8'd228, 8'd193};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd225, 8'd176, 8'd83};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd212, 8'd142, 8'd0};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd249, 8'd155, 8'd0};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd255, 8'd167, 8'd55};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd189, 8'd68, 8'd15};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd139, 8'd22, 8'd4};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd172, 8'd64, 8'd52};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd145: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd230, 8'd231, 8'd217};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd249, 8'd191, 8'd180};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd155, 8'd40, 8'd45};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd165, 8'd3, 8'd16};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd196, 8'd27, 8'd20};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd194, 8'd58, 8'd8};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd154, 8'd67};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd254, 8'd150, 8'd39};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd246, 8'd157, 8'd31};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd220, 8'd151, 8'd50};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd220, 8'd179};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd249, 8'd243, 8'd193};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd223, 8'd195, 8'd111};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd203, 8'd152, 8'd35};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd201, 8'd133, 8'd0};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd217, 8'd139, 8'd0};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd216, 8'd140, 8'd0};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd216, 8'd142, 8'd0};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd218, 8'd143, 8'd0};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd218, 8'd147, 8'd5};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd220, 8'd148, 8'd10};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd220, 8'd151, 8'd14};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd220, 8'd152, 8'd17};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd218, 8'd163, 8'd34};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd224, 8'd170, 8'd38};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd221, 8'd167, 8'd33};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd213, 8'd159, 8'd24};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd215, 8'd162, 8'd24};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd224, 8'd171, 8'd31};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd230, 8'd177, 8'd37};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd231, 8'd178, 8'd36};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd230, 8'd174, 8'd35};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd228, 8'd175, 8'd35};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd226, 8'd177, 8'd36};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd228, 8'd181, 8'd41};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd233, 8'd184, 8'd47};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd236, 8'd184, 8'd49};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd237, 8'd179, 8'd46};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd235, 8'd175, 8'd43};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd231, 8'd179, 8'd57};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd231, 8'd179, 8'd57};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd232, 8'd180, 8'd58};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd233, 8'd183, 8'd60};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd236, 8'd186, 8'd63};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd237, 8'd189, 8'd65};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd237, 8'd189, 8'd65};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd237, 8'd189, 8'd65};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd240, 8'd192, 8'd64};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd249, 8'd201, 8'd73};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd243, 8'd198, 8'd71};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd242, 8'd197, 8'd70};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd251, 8'd207, 8'd82};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd248, 8'd207, 8'd83};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd244, 8'd203, 8'd79};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd253, 8'd212, 8'd88};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd234, 8'd202, 8'd79};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd240, 8'd206, 8'd83};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd247, 8'd211, 8'd91};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd247, 8'd207, 8'd93};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd242, 8'd202, 8'd89};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd243, 8'd207, 8'd97};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd241, 8'd211, 8'd101};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd231, 8'd203, 8'd94};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd249, 8'd217, 8'd116};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd244, 8'd212, 8'd109};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd245, 8'd213, 8'd104};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd243, 8'd211, 8'd100};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd242, 8'd210, 8'd99};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd250, 8'd217, 8'd110};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd254, 8'd222, 8'd121};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd249, 8'd216, 8'd119};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd248, 8'd217, 8'd124};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd248, 8'd219, 8'd127};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd248, 8'd221, 8'd132};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd248, 8'd223, 8'd139};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd249, 8'd226, 8'd148};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd249, 8'd229, 8'd156};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd250, 8'd231, 8'd162};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd250, 8'd233, 8'd164};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd252, 8'd228, 8'd156};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd247, 8'd217, 8'd131};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd236, 8'd198, 8'd89};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd221, 8'd178, 8'd47};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd211, 8'd166, 8'd25};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd207, 8'd166, 8'd26};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd211, 8'd174, 8'd41};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd217, 8'd183, 8'd59};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd251, 8'd238, 8'd196};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd253, 8'd242, 8'd212};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd255, 8'd215, 8'd166};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd230, 8'd174, 8'd79};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd246, 8'd179, 8'd39};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd242, 8'd160, 8'd24};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd227, 8'd135, 8'd48};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd153, 8'd63, 8'd29};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd190, 8'd113, 8'd107};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd254, 8'd188, 8'd189};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd146: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd254, 8'd196, 8'd192};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd202, 8'd99, 8'd102};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd142, 8'd14, 8'd5};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd155, 8'd26, 8'd0};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd138, 8'd73};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd245, 8'd147, 8'd36};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd241, 8'd156, 8'd11};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd223, 8'd159, 8'd23};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd255, 8'd218, 8'd152};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd247, 8'd230, 8'd176};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd217, 8'd180, 8'd102};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd191, 8'd142, 8'd50};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd198, 8'd131, 8'd24};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd199, 8'd132, 8'd25};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd200, 8'd133, 8'd26};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd200, 8'd136, 8'd28};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd200, 8'd138, 8'd29};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd202, 8'd139, 8'd33};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd202, 8'd141, 8'd34};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd203, 8'd142, 8'd35};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd212, 8'd167, 8'd52};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd205, 8'd160, 8'd45};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd210, 8'd165, 8'd48};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd211, 8'd166, 8'd49};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd197, 8'd152, 8'd33};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd190, 8'd146, 8'd25};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd198, 8'd154, 8'd33};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd203, 8'd159, 8'd38};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd202, 8'd157, 8'd40};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd198, 8'd156, 8'd38};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd198, 8'd156, 8'd38};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd201, 8'd159, 8'd41};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd208, 8'd161, 8'd45};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd213, 8'd157, 8'd44};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd211, 8'd149, 8'd38};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd207, 8'd141, 8'd31};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd208, 8'd145, 8'd50};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd207, 8'd147, 8'd51};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd207, 8'd149, 8'd52};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd206, 8'd150, 8'd53};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd206, 8'd152, 8'd54};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd206, 8'd154, 8'd55};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd206, 8'd156, 8'd57};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd207, 8'd159, 8'd59};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd210, 8'd157, 8'd55};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd216, 8'd163, 8'd61};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd213, 8'd161, 8'd60};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd212, 8'd160, 8'd59};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd218, 8'd168, 8'd69};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd216, 8'd168, 8'd70};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd214, 8'd166, 8'd68};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd217, 8'd171, 8'd75};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd206, 8'd168, 8'd67};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd219, 8'd180, 8'd79};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd223, 8'd179, 8'd82};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd218, 8'd172, 8'd76};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd220, 8'd174, 8'd80};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd220, 8'd175, 8'd82};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd211, 8'd170, 8'd78};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd206, 8'd170, 8'd76};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd212, 8'd181, 8'd88};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd206, 8'd176, 8'd80};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd198, 8'd169, 8'd69};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd201, 8'd172, 8'd70};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd210, 8'd181, 8'd79};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd207, 8'd178, 8'd78};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd202, 8'd172, 8'd76};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd206, 8'd175, 8'd82};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd205, 8'd174, 8'd83};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd204, 8'd175, 8'd83};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd204, 8'd177, 8'd86};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd205, 8'd179, 8'd92};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd206, 8'd182, 8'd96};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd206, 8'd185, 8'd102};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd205, 8'd187, 8'd105};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd206, 8'd188, 8'd106};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd207, 8'd177, 8'd113};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd208, 8'd174, 8'd100};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd202, 8'd165, 8'd76};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd190, 8'd149, 8'd44};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd181, 8'd140, 8'd32};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd193, 8'd156, 8'd52};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd221, 8'd190, 8'd97};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd247, 8'd220, 8'd133};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd255, 8'd224, 8'd166};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd205, 8'd151, 8'd65};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd221, 8'd163, 8'd55};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd229, 8'd166, 8'd71};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd245, 8'd185, 8'd133};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd213, 8'd166, 8'd156};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd147: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd186, 8'd114, 8'd102};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd142, 8'd47, 8'd15};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd233, 8'd127, 8'd77};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd236, 8'd150, 8'd49};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd229, 8'd155, 8'd6};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd219, 8'd163, 8'd8};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd251, 8'd213, 8'd130};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd254, 8'd246, 8'd223};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd245, 8'd225, 8'd188};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd231, 8'd202, 8'd158};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd233, 8'd208, 8'd168};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd234, 8'd209, 8'd168};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd234, 8'd211, 8'd167};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd235, 8'd213, 8'd166};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd236, 8'd214, 8'd165};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd237, 8'd215, 8'd165};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd238, 8'd217, 8'd164};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd238, 8'd217, 8'd164};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd249, 8'd222, 8'd169};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd238, 8'd211, 8'd158};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd239, 8'd212, 8'd159};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd244, 8'd217, 8'd164};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd208, 8'd181, 8'd126};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd140, 8'd113, 8'd58};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd107, 8'd80, 8'd25};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd120, 8'd93, 8'd38};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd124, 8'd95, 8'd51};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd125, 8'd97, 8'd50};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd126, 8'd98, 8'd51};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd129, 8'd97, 8'd50};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd129, 8'd91, 8'd44};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd129, 8'd82, 8'd36};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd128, 8'd71, 8'd28};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd126, 8'd65, 8'd21};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd127, 8'd65, 8'd28};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd129, 8'd67, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd127, 8'd67, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd123, 8'd68, 8'd29};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd119, 8'd67, 8'd27};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd118, 8'd69, 8'd28};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd121, 8'd74, 8'd32};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd123, 8'd78, 8'd36};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd121, 8'd68, 8'd26};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd123, 8'd70, 8'd28};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd122, 8'd69, 8'd27};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd122, 8'd70, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd123, 8'd74, 8'd34};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd123, 8'd74, 8'd34};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd122, 8'd74, 8'd36};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd124, 8'd76, 8'd38};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd118, 8'd80, 8'd35};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd121, 8'd80, 8'd36};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd112, 8'd67, 8'd25};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd113, 8'd66, 8'd24};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd125, 8'd77, 8'd37};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd119, 8'd74, 8'd33};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd112, 8'd70, 8'd28};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd120, 8'd83, 8'd41};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd127, 8'd101, 8'd66};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd122, 8'd98, 8'd60};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd111, 8'd89, 8'd48};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd110, 8'd91, 8'd48};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd109, 8'd90, 8'd47};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd97, 8'd76, 8'd33};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd114, 8'd91, 8'd49};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd162, 8'd137, 8'd96};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd241, 8'd217, 8'd173};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd241, 8'd218, 8'd174};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd242, 8'd219, 8'd177};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd242, 8'd221, 8'd178};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd242, 8'd223, 8'd180};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd243, 8'd226, 8'd182};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd242, 8'd228, 8'd183};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd242, 8'd228, 8'd183};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd241, 8'd215, 8'd192};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd247, 8'd220, 8'd191};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd251, 8'd221, 8'd185};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd243, 8'd211, 8'd170};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd230, 8'd202, 8'd162};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd234, 8'd210, 8'd176};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd252, 8'd235, 8'd209};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd251, 8'd217, 8'd169};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd208, 8'd174, 8'd113};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd232, 8'd197, 8'd131};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd251, 8'd215, 8'd163};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd148: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd239, 8'd193, 8'd169};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd216, 8'd152, 8'd114};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd238, 8'd176, 8'd101};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd220, 8'd165, 8'd38};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd212, 8'd165, 8'd27};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd235, 8'd199, 8'd125};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd147, 8'd142, 8'd138};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd64, 8'd59, 8'd55};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd51, 8'd46, 8'd42};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd56, 8'd50, 8'd60};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd61, 8'd55, 8'd65};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd65, 8'd60, 8'd66};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd65, 8'd54, 8'd60};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd58, 8'd42, 8'd45};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd53, 8'd27, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd52, 8'd16, 8'd20};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd53, 8'd11, 8'd15};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd60, 8'd10, 8'd3};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd61, 8'd12, 8'd5};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd61, 8'd14, 8'd6};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd55, 8'd11, 8'd2};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd49, 8'd6, 8'd0};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd47, 8'd7, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd53, 8'd15, 8'd4};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd60, 8'd22, 8'd11};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd56, 8'd9, 8'd0};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd52, 8'd8, 8'd0};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd54, 8'd10, 8'd0};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd54, 8'd11, 8'd2};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd53, 8'd10, 8'd3};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd52, 8'd12, 8'd4};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd53, 8'd14, 8'd7};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd51, 8'd12, 8'd5};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd57, 8'd24, 8'd9};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd52, 8'd16, 8'd2};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd39, 8'd1, 8'd0};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd41, 8'd3, 8'd0};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd48, 8'd11, 8'd2};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd39, 8'd6, 8'd0};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd45, 8'd18, 8'd9};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd77, 8'd55, 8'd44};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd80, 8'd67, 8'd76};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd75, 8'd65, 8'd73};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd64, 8'd62, 8'd67};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd57, 8'd57, 8'd59};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd39, 8'd39, 8'd39};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd26, 8'd25, 8'd23};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd87, 8'd79, 8'd77};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd182, 8'd171, 8'd169};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd149: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd242, 8'd235, 8'd217};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd255, 8'd247, 8'd221};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd252, 8'd218, 8'd181};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd230, 8'd195, 8'd113};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd219, 8'd184, 8'd90};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd225, 8'd194, 8'd148};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd208, 8'd218, 8'd219};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd112, 8'd122, 8'd124};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd50, 8'd60, 8'd62};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd49, 8'd61, 8'd83};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd53, 8'd66, 8'd85};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd55, 8'd68, 8'd84};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd57, 8'd67, 8'd77};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd53, 8'd58, 8'd64};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd49, 8'd44, 8'd50};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd43, 8'd31, 8'd35};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd42, 8'd23, 8'd27};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd58, 8'd21, 8'd3};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd61, 8'd24, 8'd6};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd62, 8'd25, 8'd7};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd55, 8'd18, 8'd0};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd47, 8'd10, 8'd0};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd47, 8'd10, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd56, 8'd19, 8'd1};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd66, 8'd29, 8'd11};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd65, 8'd24, 8'd4};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd58, 8'd20, 8'd0};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd61, 8'd23, 8'd4};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd62, 8'd25, 8'd6};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd57, 8'd20, 8'd2};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd57, 8'd21, 8'd5};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd59, 8'd26, 8'd9};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd54, 8'd21, 8'd4};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd68, 8'd34, 8'd9};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd64, 8'd29, 8'd7};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd59, 8'd24, 8'd5};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd55, 8'd23, 8'd8};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd49, 8'd23, 8'd10};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd44, 8'd26, 8'd14};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd70, 8'd58, 8'd46};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd109, 8'd103, 8'd91};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd89, 8'd89, 8'd101};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd81, 8'd88, 8'd98};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd72, 8'd86, 8'd95};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd60, 8'd79, 8'd86};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd43, 8'd62, 8'd68};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd56, 8'd72, 8'd72};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd141, 8'd150, 8'd149};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd150: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd245, 8'd230, 8'd199};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd248, 8'd224, 8'd186};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd239, 8'd217, 8'd206};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd185, 8'd195, 8'd196};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd97, 8'd107, 8'd109};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd61, 8'd76, 8'd99};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd54, 8'd71, 8'd91};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd53, 8'd70, 8'd86};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd61, 8'd78, 8'd86};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd74, 8'd85, 8'd89};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd74, 8'd80, 8'd80};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd62, 8'd61, 8'd57};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd49, 8'd44, 8'd40};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd68, 8'd32, 8'd8};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd74, 8'd36, 8'd13};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd76, 8'd35, 8'd13};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd71, 8'd26, 8'd5};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd61, 8'd14, 8'd0};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd63, 8'd12, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd75, 8'd22, 8'd4};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd89, 8'd33, 8'd16};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd82, 8'd34, 8'd11};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd74, 8'd26, 8'd3};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd79, 8'd31, 8'd9};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd81, 8'd35, 8'd12};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd71, 8'd26, 8'd5};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd73, 8'd28, 8'd7};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd77, 8'd34, 8'd15};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd69, 8'd26, 8'd7};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd76, 8'd29, 8'd3};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd70, 8'd24, 8'd0};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd66, 8'd21, 8'd2};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd59, 8'd19, 8'd7};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd57, 8'd27, 8'd17};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd74, 8'd55, 8'd49};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd98, 8'd89, 8'd84};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd109, 8'd105, 8'd102};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd93, 8'd95, 8'd107};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd82, 8'd90, 8'd101};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd70, 8'd87, 8'd97};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd59, 8'd81, 8'd92};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd68, 8'd91, 8'd97};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd122, 8'd140, 8'd140};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd203, 8'd214, 8'd210};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd151: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd172, 8'd171, 8'd185};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd73, 8'd81, 8'd118};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd59, 8'd68, 8'd101};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd52, 8'd63, 8'd91};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd68, 8'd79, 8'd99};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd94, 8'd102, 8'd115};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd102, 8'd105, 8'd114};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd83, 8'd81, 8'd86};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd61, 8'd55, 8'd57};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd75, 8'd31, 8'd20};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd82, 8'd35, 8'd25};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd85, 8'd35, 8'd26};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd79, 8'd24, 8'd17};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd71, 8'd10, 8'd5};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd75, 8'd7, 8'd4};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd89, 8'd18, 8'd16};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd104, 8'd30, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd90, 8'd27, 8'd18};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd81, 8'd18, 8'd11};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd85, 8'd25, 8'd17};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd88, 8'd27, 8'd22};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd76, 8'd17, 8'd11};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd78, 8'd20, 8'd16};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd84, 8'd26, 8'd22};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd75, 8'd17, 8'd15};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd93, 8'd29, 8'd20};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd79, 8'd16, 8'd9};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd69, 8'd9, 8'd9};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd62, 8'd11, 8'd16};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd76, 8'd36, 8'd47};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd115, 8'd88, 8'd103};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd126, 8'd111, 8'd130};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd99, 8'd90, 8'd111};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd97, 8'd92, 8'd115};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd82, 8'd82, 8'd108};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd66, 8'd76, 8'd101};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd59, 8'd77, 8'd101};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd93, 8'd111, 8'd131};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd180, 8'd192, 8'd206};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd152: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd166, 8'd162, 8'd179};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd86, 8'd89, 8'd104};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd58, 8'd72, 8'd85};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd84, 8'd106, 8'd117};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd100, 8'd124, 8'd136};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd111, 8'd130, 8'd145};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd107, 8'd115, 8'd134};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd75, 8'd77, 8'd100};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd90, 8'd63, 8'd68};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd70, 8'd36, 8'd37};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd78, 8'd33, 8'd27};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd89, 8'd36, 8'd22};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd72, 8'd13, 8'd0};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd66, 8'd8, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd86, 8'd34, 8'd12};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd104, 8'd53, 8'd32};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd85, 8'd19, 8'd5};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd99, 8'd37, 8'd14};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd88, 8'd31, 8'd2};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd87, 8'd33, 8'd9};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd78, 8'd24, 8'd12};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd48, 8'd0, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd99, 8'd48, 8'd29};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd86, 8'd35, 8'd4};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd97, 8'd31, 8'd7};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd73, 8'd16, 8'd0};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd56, 8'd19, 8'd3};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd70, 8'd50, 8'd43};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd88, 8'd85};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd109, 8'd110, 8'd114};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd115, 8'd119, 8'd128};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd119, 8'd123, 8'd132};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd100, 8'd122, 8'd136};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd80, 8'd99, 8'd113};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd66, 8'd83, 8'd93};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd93, 8'd106, 8'd114};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd165, 8'd173, 8'd176};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd153: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd224, 8'd222, 8'd236};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd135, 8'd141, 8'd153};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd86, 8'd103, 8'd113};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd97, 8'd121, 8'd131};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd105, 8'd132, 8'd143};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd107, 8'd129, 8'd143};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd111, 8'd124, 8'd141};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd106, 8'd112, 8'd134};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd99, 8'd82, 8'd88};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd101, 8'd77, 8'd77};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd78, 8'd41, 8'd35};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd68, 8'd20, 8'd6};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd85, 8'd28, 8'd9};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd77, 8'd16, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd76, 8'd16, 8'd0};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd109, 8'd51, 8'd29};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd98, 8'd29, 8'd13};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd97, 8'd31, 8'd5};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd97, 8'd36, 8'd5};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd117, 8'd57, 8'd31};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd98, 8'd39, 8'd25};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd58, 8'd0, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd103, 8'd46, 8'd29};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd85, 8'd29, 8'd2};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd100, 8'd38, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd74, 8'd23, 8'd4};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd70, 8'd36, 8'd24};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd99, 8'd84, 8'd79};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd120, 8'd120, 8'd122};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd112, 8'd119, 8'd127};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd99, 8'd109, 8'd121};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd98, 8'd107, 8'd122};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd94, 8'd113, 8'd127};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd82, 8'd100, 8'd112};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd90, 8'd107, 8'd115};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd142, 8'd153, 8'd159};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd208, 8'd216, 8'd219};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd154: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd191, 8'd200, 8'd207};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd127, 8'd144, 8'd151};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd103, 8'd128, 8'd135};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd99, 8'd126, 8'd135};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd102, 8'd126, 8'd138};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd115, 8'd134, 8'd149};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd130, 8'd145, 8'd164};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd121, 8'd119, 8'd124};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd100, 8'd90, 8'd91};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd90, 8'd69, 8'd64};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd91, 8'd55, 8'd41};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd81, 8'd30, 8'd11};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd74, 8'd14, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd90, 8'd23, 8'd0};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd111, 8'd39, 8'd14};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd108, 8'd33, 8'd12};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd107, 8'd36, 8'd6};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd114, 8'd46, 8'd9};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd131, 8'd64, 8'd35};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd100, 8'd33, 8'd17};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd61, 8'd0, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd111, 8'd49, 8'd36};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd109, 8'd48, 8'd27};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd85, 8'd34, 8'd15};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd88, 8'd46, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd105, 8'd80, 8'd73};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd128, 8'd122, 8'd122};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd131, 8'd140, 8'd147};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd110, 8'd126, 8'd139};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd89, 8'd108, 8'd125};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd81, 8'd99, 8'd119};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd79, 8'd97, 8'd109};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd94, 8'd111, 8'd121};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd139, 8'd154, 8'd161};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd219};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd155: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd178, 8'd196, 8'd198};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd122, 8'd146, 8'd150};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd104, 8'd131, 8'd138};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd110, 8'd137, 8'd148};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd125, 8'd148, 8'd162};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd142, 8'd163, 8'd180};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd158, 8'd169, 8'd175};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd110, 8'd115, 8'd118};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd99, 8'd94, 8'd90};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd104, 8'd84, 8'd73};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd82, 8'd43, 8'd26};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd76, 8'd20, 8'd0};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd101, 8'd31, 8'd5};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd116, 8'd39, 8'd11};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd108, 8'd28, 8'd3};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd125, 8'd46, 8'd13};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd120, 8'd45, 8'd5};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd129, 8'd54, 8'd22};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd105, 8'd32, 8'd17};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd69, 8'd0, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd103, 8'd40, 8'd33};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd120, 8'd62, 8'd48};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd77, 8'd39, 8'd26};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd113, 8'd86, 8'd75};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd142, 8'd131, 8'd127};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd135, 8'd140, 8'd144};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd113, 8'd129, 8'd142};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd99, 8'd122, 8'd138};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd90, 8'd115, 8'd135};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd86, 8'd108, 8'd131};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd82, 8'd96, 8'd105};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd128, 8'd143, 8'd150};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd196, 8'd207, 8'd213};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd156: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd173, 8'd193, 8'd194};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd142, 8'd165, 8'd171};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd129, 8'd153, 8'd163};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd127, 8'd154, 8'd165};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd143, 8'd169, 8'd182};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd174, 8'd194, 8'd201};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd161, 8'd179, 8'd183};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd118, 8'd128, 8'd127};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd93, 8'd90, 8'd83};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd99, 8'd77, 8'd64};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd90, 8'd47, 8'd28};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd88, 8'd26, 8'd3};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd115, 8'd41, 8'd16};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd115, 8'd29, 8'd4};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd138, 8'd54, 8'd18};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd122, 8'd41, 8'd0};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd137, 8'd58, 8'd25};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd125, 8'd52, 8'd37};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd66, 8'd2, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd66, 8'd15, 8'd14};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd114, 8'd69, 8'd63};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd110, 8'd90, 8'd83};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd137, 8'd126, 8'd122};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd150, 8'd151, 8'd153};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd125, 8'd140, 8'd147};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd115, 8'd129};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd84, 8'd110, 8'd127};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd95, 8'd117, 8'd138};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd102, 8'd124, 8'd145};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd128, 8'd139, 8'd145};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd181, 8'd192, 8'd198};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd157: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd223, 8'd234, 8'd236};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd188, 8'd205, 8'd212};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd143, 8'd166, 8'd174};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd123, 8'd147, 8'd159};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd134, 8'd160, 8'd173};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd153, 8'd176, 8'd184};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd176, 8'd201, 8'd206};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd171, 8'd195, 8'd197};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd134, 8'd149, 8'd146};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd105, 8'd105, 8'd97};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd98, 8'd74, 8'd62};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd94, 8'd47, 8'd31};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd91, 8'd30, 8'd12};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd130, 8'd40, 8'd16};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd150, 8'd61, 8'd27};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd133, 8'd50, 8'd8};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd149, 8'd73, 8'd39};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd118, 8'd52, 8'd36};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd44, 8'd0, 8'd0};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd50, 8'd15, 8'd19};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd137, 8'd116, 8'd115};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd158, 8'd156, 8'd157};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd144, 8'd148, 8'd151};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd129, 8'd142, 8'd150};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd112, 8'd134, 8'd145};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd93, 8'd119, 8'd132};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd86, 8'd109, 8'd123};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd106, 8'd123, 8'd139};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd135, 8'd148, 8'd164};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd196, 8'd204, 8'd207};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd158: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd226, 8'd237, 8'd243};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd180, 8'd197, 8'd207};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd142, 8'd164, 8'd177};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd132, 8'd158, 8'd171};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd134, 8'd154, 8'd163};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd149, 8'd176, 8'd185};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd184, 8'd215, 8'd220};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd174, 8'd204, 8'd206};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd127, 8'd143, 8'd142};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd115, 8'd110, 8'd104};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd116, 8'd87, 8'd79};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd88, 8'd44, 8'd33};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd138, 8'd46, 8'd23};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd147, 8'd58, 8'd24};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd139, 8'd56, 8'd14};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd151, 8'd78, 8'd45};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd105, 8'd47, 8'd33};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd65, 8'd29, 8'd31};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd87, 8'd74, 8'd81};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd162, 8'd161, 8'd166};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd164, 8'd174, 8'd183};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd133, 8'd150, 8'd158};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd111, 8'd133, 8'd144};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd134, 8'd145};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd106, 8'd130, 8'd142};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd110, 8'd128, 8'd138};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd142, 8'd152, 8'd161};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd182, 8'd187, 8'd193};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd159: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd184, 8'd203, 8'd217};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd148, 8'd171, 8'd185};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd141, 8'd159, 8'd169};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd138, 8'd165, 8'd174};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd135, 8'd169, 8'd178};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd150, 8'd187, 8'd193};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd168, 8'd196, 8'd197};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd148, 8'd154, 8'd152};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd120, 8'd102, 8'd98};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd119, 8'd89, 8'd81};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd138, 8'd43, 8'd23};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd131, 8'd40, 8'd9};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd127, 8'd44, 8'd4};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd145, 8'd74, 8'd42};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd113, 8'd64, 8'd50};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd127, 8'd101, 8'd104};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd143, 8'd142, 8'd150};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd149, 8'd164, 8'd171};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd135, 8'd155, 8'd166};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd122, 8'd144, 8'd157};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd110, 8'd138, 8'd150};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd106, 8'd134, 8'd145};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd111, 8'd135, 8'd145};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd135, 8'd150, 8'd157};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd181, 8'd186, 8'd190};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd224, 8'd222, 8'd225};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd160: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd145, 8'd178, 8'd183};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd140, 8'd173, 8'd182};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd127, 8'd156, 8'd174};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd121, 8'd148, 8'd169};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd142, 8'd165, 8'd183};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd159, 8'd182, 8'd190};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd138, 8'd160, 8'd157};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd99, 8'd123, 8'd110};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd106, 8'd82, 8'd58};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd108, 8'd67, 8'd49};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd103, 8'd49, 8'd37};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd127, 8'd77, 8'd70};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd152, 8'd121, 8'd118};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd159, 8'd150, 8'd153};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd159, 8'd163, 8'd175};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd141, 8'd148, 8'd167};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd93, 8'd125, 8'd136};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd84, 8'd114, 8'd124};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd76, 8'd100, 8'd110};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd107, 8'd126, 8'd133};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd147, 8'd160, 8'd166};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd183, 8'd191, 8'd194};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd161: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd184, 8'd212, 8'd213};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd164, 8'd191, 8'd198};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd125, 8'd151, 8'd166};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd97, 8'd119, 8'd140};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd108, 8'd131, 8'd149};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd143, 8'd167, 8'd177};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd158, 8'd184, 8'd183};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd150, 8'd176, 8'd167};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd124, 8'd126, 8'd105};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd119, 8'd103, 8'd88};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd120, 8'd90, 8'd80};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd159, 8'd130, 8'd124};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd173, 8'd162, 8'd158};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd143, 8'd153, 8'd154};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd114, 8'd133, 8'd140};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd88, 8'd107, 8'd122};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd88, 8'd118, 8'd128};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd99, 8'd128, 8'd136};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd104, 8'd127, 8'd135};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd133, 8'd150, 8'd157};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd177, 8'd188, 8'd194};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd217, 8'd222, 8'd226};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd162: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd196, 8'd214, 8'd216};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd153, 8'd171, 8'd181};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd112, 8'd131, 8'd146};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd109, 8'd130, 8'd147};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd140, 8'd167, 8'd178};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd172, 8'd200, 8'd203};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd183, 8'd213, 8'd211};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd132, 8'd162, 8'd150};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd119, 8'd132, 8'd125};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd121, 8'd117, 8'd116};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd164, 8'd160, 8'd161};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd169, 8'd181, 8'd181};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd123, 8'd151, 8'd152};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd97, 8'd130, 8'd135};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd84, 8'd117, 8'd126};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd62, 8'd89, 8'd96};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd91, 8'd116, 8'd121};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd118, 8'd139, 8'd144};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd165, 8'd180, 8'd185};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd211, 8'd222, 8'd226};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd163: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd202, 8'd213, 8'd217};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd164, 8'd178, 8'd189};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd143, 8'd162, 8'd176};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd152, 8'd176, 8'd188};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd169, 8'd198, 8'd204};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd179, 8'd210, 8'd213};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd174, 8'd216, 8'd215};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd170, 8'd195, 8'd200};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd166, 8'd176, 8'd185};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd176, 8'd185, 8'd194};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd146, 8'd166, 8'd173};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd93, 8'd124, 8'd129};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd85, 8'd118, 8'd125};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd96, 8'd126, 8'd134};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd105, 8'd126, 8'd131};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd130, 8'd151, 8'd154};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd165, 8'd183, 8'd187};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd219, 8'd233, 8'd236};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd164: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd205, 8'd216, 8'd222};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd174, 8'd191, 8'd199};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd160, 8'd183, 8'd191};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd160, 8'd187, 8'd196};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd162, 8'd191, 8'd199};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd192, 8'd231, 8'd238};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd141, 8'd157, 8'd172};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd83, 8'd107, 8'd117};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd93, 8'd116, 8'd124};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd116, 8'd133, 8'd141};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd150, 8'd168, 8'd168};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd179, 8'd195, 8'd195};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd210, 8'd224, 8'd224};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd165: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd205, 8'd219, 8'd222};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd178, 8'd197, 8'd203};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd158, 8'd181, 8'd187};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd148, 8'd173, 8'd180};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd165, 8'd194, 8'd200};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd135, 8'd147, 8'd163};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd95, 8'd113, 8'd125};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd128, 8'd143, 8'd150};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd161, 8'd168, 8'd176};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd181, 8'd193, 8'd189};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd166: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd210, 8'd224, 8'd225};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd182, 8'd197, 8'd202};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd162, 8'd179, 8'd186};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd160, 8'd186, 8'd185};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd140, 8'd154, 8'd167};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd117, 8'd137, 8'd144};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd161, 8'd176, 8'd181};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd196, 8'd204, 8'd207};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd167: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd213, 8'd224, 8'd226};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd195, 8'd209, 8'd212};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd163, 8'd190, 8'd181};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd169, 8'd189, 8'd198};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd155, 8'd183, 8'd186};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd196, 8'd217, 8'd218};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd168: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd169: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd170: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd171: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd172: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd173: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd174: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd175: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd176: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd177: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd178: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd179: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd180: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd181: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
				`ybit'd182: begin
					case(X)
						`xbit'd0: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd1: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd2: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd3: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd4: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd5: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd6: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd7: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd8: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd9: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd10: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd11: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd12: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd13: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd14: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd15: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd16: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd17: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd18: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd19: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd20: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd21: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd22: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd23: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd24: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd25: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd26: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd27: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd28: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd29: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd30: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd31: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd32: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd33: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd34: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd35: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd36: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd37: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd38: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd39: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd40: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd41: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd42: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd43: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd44: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd45: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd46: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd47: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd48: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd49: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd50: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd51: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd52: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd53: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd54: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd55: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd56: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd57: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd58: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd59: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd60: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd61: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd62: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd63: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd64: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd65: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd66: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd67: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd68: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd69: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd70: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd71: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd72: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd73: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd74: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd75: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd76: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd77: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd78: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd79: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd80: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd81: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd82: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd83: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd84: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd85: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd86: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd87: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd88: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd89: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd90: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd91: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd92: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd93: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd94: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd95: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd96: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd97: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd98: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd99: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd100: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd101: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd102: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd103: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd104: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd105: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd106: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd107: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd108: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd109: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd110: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd111: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd112: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd113: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd114: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd115: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd116: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd117: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd118: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd119: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd120: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd121: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd122: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd123: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd124: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd125: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd126: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd127: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd128: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd129: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd130: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd131: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd132: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd133: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd134: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd135: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd136: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd137: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd138: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd139: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd140: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd141: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd142: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd143: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd144: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd145: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd146: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd147: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd148: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd149: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd150: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd151: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd152: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd153: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd154: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd155: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd156: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd157: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd158: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd159: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd160: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd161: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd162: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd163: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd164: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd165: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd166: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd167: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd168: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd169: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd170: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd171: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd172: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd173: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd174: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd175: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd176: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd177: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd178: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd179: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd180: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd181: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd182: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd183: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd184: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd185: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd186: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd187: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd188: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd189: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd190: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd191: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd192: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd193: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd194: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd195: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd196: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd197: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd198: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd199: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd200: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd201: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd202: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd203: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd204: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd205: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd206: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd207: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd208: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd209: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd210: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd211: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd212: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd213: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd214: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd215: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd216: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd217: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd218: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd219: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd220: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd221: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd222: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd223: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd224: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd225: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd226: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd227: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd228: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd229: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd230: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd231: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd232: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd233: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd234: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd235: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd236: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd237: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd238: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd239: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd240: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd241: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd242: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd243: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd244: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd245: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd246: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd247: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd248: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd249: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd250: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd251: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd252: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd253: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd254: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd255: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd256: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd257: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd258: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd259: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd260: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd261: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd262: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd263: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd264: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd265: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd266: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd267: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd268: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd269: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd270: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd271: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd272: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd273: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
						`xbit'd274: {mapR, mapG, mapB} <= {8'd19, 8'd236, 8'd30};
					endcase
				end
			endcase
		end
	end

endmodule